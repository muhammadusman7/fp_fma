// Title: Leading One Detector V 1.0 (No Changelog)
// Created: Septmeber 11, 2021
// Updated: 
//---------------------------------------------------------------------------
// This is a Verilog file that define a Leading one Detection
// 
//
//---------------------------------------------------------------------------
module lod (
    input   [105:0] in,
    output reg [6:0] lo_posdp,
    output reg [6:0] lo_possp0,
    output reg [6:0] lo_possp1,
    output reg [6:0] lo_poshp0,
    output reg [6:0] lo_poshp1,
    output reg [6:0] lo_poshp2,
    output reg [6:0] lo_poshp3
);

    reg [6:0] lo_pos0, lo_pos1, lo_pos2, lo_pos3;
    // Detect Leading one from LtR
    always @(in) begin
        // First 22:0 
        casez(in[21:0])
            22'b0_0000_0000_0000_0000_0000_1: begin lo_pos0 = 7'd105; end
            22'b0_0000_0000_0000_0000_0001_?: begin lo_pos0 = 7'd104; end
            22'b0_0000_0000_0000_0000_001?_?: begin lo_pos0 = 7'd103; end
            22'b0_0000_0000_0000_0000_01??_?: begin lo_pos0 = 7'd102; end
            22'b0_0000_0000_0000_0000_1???_?: begin lo_pos0 = 7'd101; end
            22'b0_0000_0000_0000_0001_????_?: begin lo_pos0 = 7'd100; end
            22'b0_0000_0000_0000_001?_????_?: begin lo_pos0 = 7'd99;  end
            22'b0_0000_0000_0000_01??_????_?: begin lo_pos0 = 7'd98;  end
            22'b0_0000_0000_0000_1???_????_?: begin lo_pos0 = 7'd97;  end
            22'b0_0000_0000_0001_????_????_?: begin lo_pos0 = 7'd96;  end
            22'b0_0000_0000_001?_????_????_?: begin lo_pos0 = 7'd95;  end
            22'b0_0000_0000_01??_????_????_?: begin lo_pos0 = 7'd94;  end
            22'b0_0000_0000_1???_????_????_?: begin lo_pos0 = 7'd93;  end
            22'b0_0000_0001_????_????_????_?: begin lo_pos0 = 7'd92;  end
            22'b0_0000_001?_????_????_????_?: begin lo_pos0 = 7'd91;  end
            22'b0_0000_01??_????_????_????_?: begin lo_pos0 = 7'd90;  end
            22'b0_0000_1???_????_????_????_?: begin lo_pos0 = 7'd89;  end
            22'b0_0001_????_????_????_????_?: begin lo_pos0 = 7'd88;  end
            22'b0_001?_????_????_????_????_?: begin lo_pos0 = 7'd87;  end
            22'b0_01??_????_????_????_????_?: begin lo_pos0 = 7'd86;  end
            22'b0_1???_????_????_????_????_?: begin lo_pos0 = 7'd85;  end
            22'b1_????_????_????_????_????_?: begin lo_pos0 = 7'd84;  end
            default: begin lo_pos0 = 7'd127; end
        endcase
        if(lo_pos0 == 7'd127) begin
            lo_poshp0 = lo_pos0;
        end else begin
            lo_poshp0 = lo_pos0 + 7'b0101100;   // 2'comp of 84
        end
        
        // Second 50:23 
        casez(in[49:22])
            28'b0_0000_0000_0000_0000_0000_0000_001: begin lo_pos1 = 7'd83; end
            28'b0_0000_0000_0000_0000_0000_0000_01?: begin lo_pos1 = 7'd82; end
            28'b0_0000_0000_0000_0000_0000_0000_1??: begin lo_pos1 = 7'd81; end
            28'b0_0000_0000_0000_0000_0000_0001_???: begin lo_pos1 = 7'd80; end
            28'b0_0000_0000_0000_0000_0000_001?_???: begin lo_pos1 = 7'd79; end
            28'b0_0000_0000_0000_0000_0000_01??_???: begin lo_pos1 = 7'd78; end
            28'b0_0000_0000_0000_0000_0000_1???_???: begin lo_pos1 = 7'd77; end
            28'b0_0000_0000_0000_0000_0001_????_???: begin lo_pos1 = 7'd76; end
            28'b0_0000_0000_0000_0000_001?_????_???: begin lo_pos1 = 7'd75; end
            28'b0_0000_0000_0000_0000_01??_????_???: begin lo_pos1 = 7'd74; end
            28'b0_0000_0000_0000_0000_1???_????_???: begin lo_pos1 = 7'd73; end
            28'b0_0000_0000_0000_0001_????_????_???: begin lo_pos1 = 7'd72; end
            28'b0_0000_0000_0000_001?_????_????_???: begin lo_pos1 = 7'd71;  end
            28'b0_0000_0000_0000_01??_????_????_???: begin lo_pos1 = 7'd70;  end
            28'b0_0000_0000_0000_1???_????_????_???: begin lo_pos1 = 7'd69;  end
            28'b0_0000_0000_0001_????_????_????_???: begin lo_pos1 = 7'd68;  end
            28'b0_0000_0000_001?_????_????_????_???: begin lo_pos1 = 7'd67;  end
            28'b0_0000_0000_01??_????_????_????_???: begin lo_pos1 = 7'd66;  end
            28'b0_0000_0000_1???_????_????_????_???: begin lo_pos1 = 7'd65;  end
            28'b0_0000_0001_????_????_????_????_???: begin lo_pos1 = 7'd64;  end
            28'b0_0000_001?_????_????_????_????_???: begin lo_pos1 = 7'd63;  end
            28'b0_0000_01??_????_????_????_????_???: begin lo_pos1 = 7'd62;  end
            28'b0_0000_1???_????_????_????_????_???: begin lo_pos1 = 7'd61;  end
            28'b0_0001_????_????_????_????_????_???: begin lo_pos1 = 7'd60;  end
            28'b0_001?_????_????_????_????_????_???: begin lo_pos1 = 7'd59;  end
            28'b0_01??_????_????_????_????_????_???: begin lo_pos1 = 7'd58;  end
            28'b0_1???_????_????_????_????_????_???: begin lo_pos1 = 7'd57;  end
            28'b1_????_????_????_????_????_????_???: begin lo_pos1 = 7'd56;  end
            default: begin lo_pos1 = 7'd127; end
        endcase
        if(lo_pos1 == 7'd127) begin
            lo_poshp1 = lo_pos1;
        end else begin
            lo_poshp1 = lo_pos1 + 7'b1001000;   // 2'comp of 56
        end

        if( lo_pos1 < lo_pos0) begin
            lo_possp0 = lo_pos1 + 7'b1000110;      // 2'comp of 58
        end else if (lo_pos0 == 7'd127) begin
            lo_possp0 = lo_pos0;
        end else begin
            lo_possp0 = lo_pos0 + 7'b1000110;
        end

        // Third 78:51
        casez(in[77:50])
            28'b0_0000_0000_0000_0000_0000_0000_001: begin lo_pos2 = 7'd55; end
            28'b0_0000_0000_0000_0000_0000_0000_01?: begin lo_pos2 = 7'd54; end
            28'b0_0000_0000_0000_0000_0000_0000_1??: begin lo_pos2 = 7'd53; end
            28'b0_0000_0000_0000_0000_0000_0001_???: begin lo_pos2 = 7'd52; end
            28'b0_0000_0000_0000_0000_0000_001?_???: begin lo_pos2 = 7'd51; end
            28'b0_0000_0000_0000_0000_0000_01??_???: begin lo_pos2 = 7'd50; end
            28'b0_0000_0000_0000_0000_0000_1???_???: begin lo_pos2 = 7'd49; end
            28'b0_0000_0000_0000_0000_0001_????_???: begin lo_pos2 = 7'd48; end
            28'b0_0000_0000_0000_0000_001?_????_???: begin lo_pos2 = 7'd47; end
            28'b0_0000_0000_0000_0000_01??_????_???: begin lo_pos2 = 7'd46; end
            28'b0_0000_0000_0000_0000_1???_????_???: begin lo_pos2 = 7'd45; end
            28'b0_0000_0000_0000_0001_????_????_???: begin lo_pos2 = 7'd44; end
            28'b0_0000_0000_0000_001?_????_????_???: begin lo_pos2 = 7'd43; end
            28'b0_0000_0000_0000_01??_????_????_???: begin lo_pos2 = 7'd42; end
            28'b0_0000_0000_0000_1???_????_????_???: begin lo_pos2 = 7'd41; end
            28'b0_0000_0000_0001_????_????_????_???: begin lo_pos2 = 7'd40; end
            28'b0_0000_0000_001?_????_????_????_???: begin lo_pos2 = 7'd39; end
            28'b0_0000_0000_01??_????_????_????_???: begin lo_pos2 = 7'd38; end
            28'b0_0000_0000_1???_????_????_????_???: begin lo_pos2 = 7'd37; end
            28'b0_0000_0001_????_????_????_????_???: begin lo_pos2 = 7'd36; end
            28'b0_0000_001?_????_????_????_????_???: begin lo_pos2 = 7'd35; end
            28'b0_0000_01??_????_????_????_????_???: begin lo_pos2 = 7'd34; end
            28'b0_0000_1???_????_????_????_????_???: begin lo_pos2 = 7'd33; end
            28'b0_0001_????_????_????_????_????_???: begin lo_pos2 = 7'd32; end
            28'b0_001?_????_????_????_????_????_???: begin lo_pos2 = 7'd31; end
            28'b0_01??_????_????_????_????_????_???: begin lo_pos2 = 7'd30; end
            28'b0_1???_????_????_????_????_????_???: begin lo_pos2 = 7'd29; end
            28'b1_????_????_????_????_????_????_???: begin lo_pos2 = 7'd28; end
            default: begin lo_pos2 = 7'd127; end
        endcase
        if(lo_pos2 == 7'd127) begin
            lo_poshp2 = lo_pos2;
        end else begin
            lo_poshp2 = lo_pos2 + 7'b1100100;   // 2'comp of 28
        end

        // Fourth 106:79
        casez(in[105:78])
            28'b0_0000_0000_0000_0000_0000_0000_001: begin lo_pos3 = 7'd27; end
            28'b0_0000_0000_0000_0000_0000_0000_01?: begin lo_pos3 = 7'd26; end
            28'b0_0000_0000_0000_0000_0000_0000_1??: begin lo_pos3 = 7'd25; end
            28'b0_0000_0000_0000_0000_0000_0001_???: begin lo_pos3 = 7'd24; end
            28'b0_0000_0000_0000_0000_0000_001?_???: begin lo_pos3 = 7'd23; end
            28'b0_0000_0000_0000_0000_0000_01??_???: begin lo_pos3 = 7'd22; end
            28'b0_0000_0000_0000_0000_0000_1???_???: begin lo_pos3 = 7'd21; end
            28'b0_0000_0000_0000_0000_0001_????_???: begin lo_pos3 = 7'd20; end
            28'b0_0000_0000_0000_0000_001?_????_???: begin lo_pos3 = 7'd19; end
            28'b0_0000_0000_0000_0000_01??_????_???: begin lo_pos3 = 7'd18; end
            28'b0_0000_0000_0000_0000_1???_????_???: begin lo_pos3 = 7'd17; end
            28'b0_0000_0000_0000_0001_????_????_???: begin lo_pos3 = 7'd16; end
            28'b0_0000_0000_0000_001?_????_????_???: begin lo_pos3 = 7'd15; end
            28'b0_0000_0000_0000_01??_????_????_???: begin lo_pos3 = 7'd14; end
            28'b0_0000_0000_0000_1???_????_????_???: begin lo_pos3 = 7'd13; end
            28'b0_0000_0000_0001_????_????_????_???: begin lo_pos3 = 7'd12; end
            28'b0_0000_0000_001?_????_????_????_???: begin lo_pos3 = 7'd11; end
            28'b0_0000_0000_01??_????_????_????_???: begin lo_pos3 = 7'd10; end
            28'b0_0000_0000_1???_????_????_????_???: begin lo_pos3 = 7'd9;  end
            28'b0_0000_0001_????_????_????_????_???: begin lo_pos3 = 7'd8;  end
            28'b0_0000_001?_????_????_????_????_???: begin lo_pos3 = 7'd7;  end
            28'b0_0000_01??_????_????_????_????_???: begin lo_pos3 = 7'd6;  end
            28'b0_0000_1???_????_????_????_????_???: begin lo_pos3 = 7'd5;  end
            28'b0_0001_????_????_????_????_????_???: begin lo_pos3 = 7'd4;  end
            28'b0_001?_????_????_????_????_????_???: begin lo_pos3 = 7'd3;  end
            28'b0_01??_????_????_????_????_????_???: begin lo_pos3 = 7'd2;  end
            28'b0_1???_????_????_????_????_????_???: begin lo_pos3 = 7'd1;  end
            28'b1_????_????_????_????_????_????_???: begin lo_pos3 = 7'd0;  end
            default: begin lo_pos3 = 7'd127; end
        endcase
        lo_poshp3 = lo_pos3;
        if(lo_pos3 < lo_pos2) begin
            lo_possp1 = lo_pos3;
            lo_posdp  = lo_pos3;
        end else if(lo_pos2 < lo_pos1) begin
            lo_posdp  = lo_pos2;
            lo_possp1 = lo_pos2;
        end else if(lo_pos1 < lo_pos0) begin
            lo_posdp  = lo_pos1;
            lo_possp1 = lo_pos2;
        end else begin
            lo_posdp  = lo_pos0;
            lo_possp1 = lo_pos2;
        end
    end

endmodule