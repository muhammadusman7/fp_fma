// Title: Booth 53 Multiplier (No Changelog)
// Created: Septmeber 11, 2021
// Updated: 
//---------------------------------------------------------------------------
// This is a Verilog file that define a Modified Booth Multiplication for radix-4
// partial product are compressed with Wallace tree reduction
//
//---------------------------------------------------------------------------
module multiplier53Booth #(parameter WIDTH = 53) (
    input       [WIDTH-1:0]     multiplicand,
    input       [WIDTH-1:0]     multiplier,
    input       [1:0]           mode,
    output reg  [2*WIDTH-1:0]   p0, p1
);

    wire [WIDTH:0] pp_in, pp_n, pp_2, pp_2n, pp_zero;
    wire [WIDTH/2:0] comp;
    wire [WIDTH+1:0] temp_multiplier;
    wire [WIDTH:0]   pp  [WIDTH/2:0];
    reg [WIDTH:0]   p  [WIDTH/2:0];

    assign temp_multiplier = {1'b0, multiplier, 1'b0};

    // Get basic partial products
    boothPP #(.WIDTH(WIDTH)) bPP (
        .in(multiplicand), .out_in(pp_in), .out_in_n(pp_n), .out_in_2(pp_2),
        .out_in_2n(pp_2n), .out_zero(pp_zero) );

    // Get partial produts for each row
    genvar i;
    generate
        for (i=0; i <= WIDTH/2; i = i+1) begin
            boothPPCal #(.WIDTH(WIDTH)) pp (.pp(pp_in), .pp_n(pp_n), .pp_2(pp_2), .pp_2n(pp_2n),
                .pp_zero(pp_zero), .booth({temp_multiplier[2*(i+1)], temp_multiplier[2*(i+1)-1], 
                temp_multiplier[2*(i+1)-2]}), .comp(comp[i]), .out(pp[i]) );
        end
    endgenerate
    
    wire [1462:0] s, c;

    always @(*) begin

        if(mode == 2'b01) begin
            p[26] = {pp[26][53:42], 42'b0};
            p[25] = {pp[25][53:42], 42'b0};
            p[24] = {pp[24][53:42], 42'b0};
            p[23] = {pp[23][53:42], 42'b0};
            p[22] = {pp[22][53:42], 42'b0};
            p[21] = {pp[21][53:42], 42'b0};
            p[20] = pp[20];
            p[19] = {14'b0, pp[19][39:28], 28'b0};
            p[18] = {14'b0, pp[18][39:28], 28'b0};
            p[17] = {14'b0, pp[17][39:28], 28'b0};
            p[16] = {14'b0, pp[16][39:28], 28'b0};
            p[15] = {14'b0, pp[15][39:28], 28'b0};
            p[14] = {14'b0, pp[14][39:28], 28'b0};
            p[13] = pp[13];
            p[12] = {28'b0, pp[12][25:14], 14'b0};
            p[11] = {28'b0, pp[11][25:14], 14'b0};
            p[10] = {28'b0, pp[10][25:14], 14'b0};
            p[9] = {28'b0, pp[9][25:14], 14'b0};
            p[8] = {28'b0, pp[8][25:14], 14'b0};
            p[7] = {28'b0, pp[7][25:14], 14'b0};
            p[6] = pp[6];
            p[5] = {42'b0, pp[5][11:0]};
            p[4] = {42'b0, pp[4][11:0]};
            p[3] = {42'b0, pp[3][11:0]};
            p[2] = {42'b0, pp[2][11:0]};
            p[1] = {42'b0, pp[1][11:0]};
            p[0] = {42'b0, pp[0][11:0]};
        end

        else if(mode == 2'b10) begin
            p[12] = {29'b0, pp[12][24:0]};
            p[11] = {29'b0, pp[11][24:0]};
            p[10] = {29'b0, pp[10][24:0]};
            p[9] = {29'b0, pp[9][24:0]};
            p[8] = {29'b0, pp[8][24:0]};
            p[7] = {29'b0, pp[7][24:0]};
            p[6] = {29'b0, pp[6][24:0]};
            p[5] = {29'b0, pp[5][24:0]};
            p[4] = {29'b0, pp[4][24:0]};
            p[3] = {29'b0, pp[3][24:0]};
            p[2] = {29'b0, pp[2][24:0]};
            p[1] = {29'b0, pp[1][24:0]};
            p[0] = {29'b0, pp[0][24:0]};
            p[13] = pp[13];
            p[26] = {pp[26][53:29], 29'b0};
            p[25] = {pp[25][53:29], 29'b0};
            p[24] = {pp[24][53:29], 29'b0};
            p[23] = {pp[23][53:29], 29'b0};
            p[22] = {pp[22][53:29], 29'b0};
            p[21] = {pp[21][53:29], 29'b0};
            p[20] = {pp[20][53:29], 29'b0};
            p[19] = {pp[19][53:29], 29'b0};
            p[18] = {pp[18][53:29], 29'b0};
            p[17] = {pp[17][53:29], 29'b0};
            p[16] = {pp[16][53:29], 29'b0};
            p[15] = {pp[15][53:29], 29'b0};
            p[14] = {pp[14][53:29], 29'b0};
        end
        else begin
            p[0][53:0] = pp[0][53:0];
            p[1][53:0] = pp[1][53:0];
            p[2][53:0] = pp[2][53:0];
            p[3][53:0] = pp[3][53:0];
            p[4][53:0] = pp[4][53:0];
            p[5][53:0] = pp[5][53:0];
            p[6][53:0] = pp[6][53:0];
            p[7][53:0] = pp[7][53:0];
            p[8][53:0] = pp[8][53:0];
            p[9][53:0] = pp[9][53:0];
            p[10][53:0] = pp[10][53:0];
            p[11][53:0] = pp[11][53:0];
            p[12][53:0] = pp[12][53:0];
            p[13][53:0] = pp[13][53:0];
            p[14][53:0] = pp[14][53:0];
            p[15][53:0] = pp[15][53:0];
            p[16][53:0] = pp[16][53:0];
            p[17][53:0] = pp[17][53:0];
            p[18][53:0] = pp[18][53:0];
            p[19][53:0] = pp[19][53:0];
            p[20][53:0] = pp[20][53:0];
            p[21][53:0] = pp[21][53:0];
            p[22][53:0] = pp[22][53:0];
            p[23][53:0] = pp[23][53:0];
            p[24][53:0] = pp[24][53:0];
            p[25][53:0] = pp[25][53:0];
            p[26][53:0] = pp[26][53:0];
        end

            p0 = {s[1094], s[855], s[1232], s[1093], s[1231], s[1462], s[1461], s[1401], s[1342], s[1460], s[1459], s[1458], s[1457], s[1456], s[1400], s[1455], s[1454], s[1453], s[1452], s[1451], s[1450], s[1449], s[1448], s[1447], s[1446], s[1445], s[1444], s[1443], s[1442], s[1441], s[1440], s[1439], s[1438], s[1437], s[1436], s[1435], s[1434], s[1433], s[1432], s[1431], s[1430], s[1429], s[1428], s[1427], s[1426], s[1425], s[1424], s[1423], s[1422], s[1421], s[1420], s[1419], s[1418], s[1417], s[1416], s[1415], s[1414], s[1413], s[1412], s[1411], s[1410], s[1409], s[1408], s[1407], s[1406], s[1405], s[1404], s[1355], s[1354], s[1353], s[1352], s[1351], s[1350], s[1349], s[1348], s[1403], s[1347], s[1346], s[1345], s[1402], s[1344], s[1240], s[1239], s[1238], s[1237], s[1236], s[1235], s[1343], s[1234], s[1101], s[1100], s[1099], s[1098], s[1233], s[1097], s[859], s[858], s[1096], s[857], s[510], s[1095], s[856], s[509], s[0], p[00][01], p[00][00]};
            p1 = {1'b0, c[1232], 1'b0, c[1231], c[1462], c[1461], 1'b0, 1'b0, c[1460], c[1459], c[1458], c[1457], c[1456], 1'b0, c[1455], c[1454], c[1453], c[1452], c[1451], c[1450], c[1449], c[1448], c[1447], c[1446], c[1445], c[1444], c[1443], c[1442], c[1441], c[1440], c[1439], c[1438], c[1437], c[1436], c[1435], c[1434], c[1433], c[1432], c[1431], c[1430], c[1429], c[1428], c[1427], c[1426], c[1425], c[1424], c[1423], c[1422], c[1421], c[1420], c[1419], c[1418], c[1417], c[1416], c[1415], c[1414], c[1413], c[1412], c[1411], c[1410], c[1409], c[1408], c[1407], c[1406], c[1405], c[1404], 1'b0, c[1354], c[1353], c[1352], c[1351], c[1350], c[1349], c[1348], c[1403], 1'b0, c[1346], c[1345], c[1402], 1'b0, 1'b0, c[1239], c[1238], c[1237], c[1236], c[1235], c[1343], 1'b0, 1'b0, c[1100], c[1099], c[1098], c[1233], 1'b0, 1'b0, c[858], c[1096], 1'b0, 1'b0, c[1095], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, comp[0]};
    
    end



    // Wallace tree reduction
    // Stage 1 Reduction
    fullAdder fa1 (.a(p[00][02]), .b(p[01][00]), .c_in(comp[1]), .s(s[0]), .c_out(c[0]));
    fullAdder fa2 (.a(p[00][04]), .b(p[01][02]), .c_in(p[02][00]), .s(s[1]), .c_out(c[1]));
    fullAdder fa3 (.a(p[00][05]), .b(p[01][03]), .c_in(p[02][01]), .s(s[2]), .c_out(c[2]));
    fullAdder fa4 (.a(p[00][06]), .b(p[01][04]), .c_in(p[02][02]), .s(s[3]), .c_out(c[3]));
    halfAdder ha1 (.a(p[03][00]), .b(comp[3]), .s(s[4]), .c_out(c[4]));
    fullAdder fa5 (.a(p[00][07]), .b(p[01][05]), .c_in(p[02][03]), .s(s[5]), .c_out(c[5]));
    fullAdder fa6 (.a(p[00][08]), .b(p[01][06]), .c_in(p[02][04]), .s(s[6]), .c_out(c[6]));
    fullAdder fa7 (.a(p[03][02]), .b(p[04][00]), .c_in(comp[4]), .s(s[7]), .c_out(c[7]));
    fullAdder fa8 (.a(p[00][09]), .b(p[01][07]), .c_in(p[02][05]), .s(s[8]), .c_out(c[8]));
    halfAdder ha2 (.a(p[03][03]), .b(p[04][01]), .s(s[9]), .c_out(c[9]));
    fullAdder fa9 (.a(p[00][10]), .b(p[01][08]), .c_in(p[02][06]), .s(s[10]), .c_out(c[10]));
    fullAdder fa10 (.a(p[03][04]), .b(p[04][02]), .c_in(p[05][00]), .s(s[11]), .c_out(c[11]));
    fullAdder fa11 (.a(p[00][11]), .b(p[01][09]), .c_in(p[02][07]), .s(s[12]), .c_out(c[12]));
    fullAdder fa12 (.a(p[03][05]), .b(p[04][03]), .c_in(p[05][01]), .s(s[13]), .c_out(c[13]));
    fullAdder fa13 (.a(mode == 2'b01 ? comp[0] : p[00][12]), .b(p[01][10]), .c_in(p[02][08]), .s(s[14]), .c_out(c[14]));
    fullAdder fa14 (.a(p[03][06]), .b(p[04][04]), .c_in(p[05][02]), .s(s[15]), .c_out(c[15]));
    halfAdder ha3 (.a(p[06][00]), .b(mode == 2'b01 ? 1'b0 : comp[6]), .s(s[16]), .c_out(c[16]));
    fullAdder fa15 (.a(mode == 2'b01 ? comp[0] : p[00][13]), .b(p[01][11]), .c_in(p[02][09]), .s(s[17]), .c_out(c[17]));
    fullAdder fa16 (.a(p[03][07]), .b(p[04][05]), .c_in(p[05][03]), .s(s[18]), .c_out(c[18]));
    fullAdder fa17 (.a(mode == 2'b01 ? ~comp[0] : p[00][14]), .b(mode == 2'b01 ? ~comp[1] : p[01][12]), .c_in(p[02][10]), .s(s[19]), .c_out(c[19]));
    fullAdder fa18 (.a(p[03][08]), .b(p[04][06]), .c_in(p[05][04]), .s(s[20]), .c_out(c[20]));
    fullAdder fa19 (.a(p[06][02]), .b(p[07][00]), .c_in(mode == 2'b01 ? 1'b0 : comp[7]), .s(s[21]), .c_out(c[21]));
    fullAdder fa20 (.a(p[00][15]), .b(mode == 2'b01 ? 1'b1 : p[01][13]), .c_in(p[02][11]), .s(s[22]), .c_out(c[22]));
    fullAdder fa21 (.a(p[03][09]), .b(p[04][07]), .c_in(p[05][05]), .s(s[23]), .c_out(c[23]));
    halfAdder ha4 (.a(p[06][03]), .b(p[07][01]), .s(s[24]), .c_out(c[24]));
    fullAdder fa22 (.a(p[00][16]), .b(p[01][14]), .c_in(mode == 2'b01 ? ~comp[2] : p[02][12]), .s(s[25]), .c_out(c[25]));
    fullAdder fa23 (.a(p[03][10]), .b(p[04][08]), .c_in(p[05][06]), .s(s[26]), .c_out(c[26]));
    fullAdder fa24 (.a(p[06][04]), .b(p[07][02]), .c_in(p[08][00]), .s(s[27]), .c_out(c[27]));
    fullAdder fa25 (.a(p[00][17]), .b(p[01][15]), .c_in(mode == 2'b01 ? 1'b1 : p[02][13]), .s(s[28]), .c_out(c[28]));
    fullAdder fa26 (.a(p[03][11]), .b(p[04][09]), .c_in(p[05][07]), .s(s[29]), .c_out(c[29]));
    fullAdder fa27 (.a(p[06][05]), .b(p[07][03]), .c_in(p[08][01]), .s(s[30]), .c_out(c[30]));
    fullAdder fa28 (.a(p[00][18]), .b(p[01][16]), .c_in(p[02][14]), .s(s[31]), .c_out(c[31]));
    fullAdder fa29 (.a(mode == 2'b01 ? ~comp[3] : p[03][12]), .b(p[04][10]), .c_in(p[05][08]), .s(s[32]), .c_out(c[32]));
    fullAdder fa30 (.a(p[06][06]), .b(p[07][04]), .c_in(p[08][02]), .s(s[33]), .c_out(c[33]));
    halfAdder ha5 (.a(p[09][00]), .b(mode == 2'b01 ? 1'b0 : comp[9]), .s(s[34]), .c_out(c[34]));
    fullAdder fa31 (.a(p[00][19]), .b(p[01][17]), .c_in(p[02][15]), .s(s[35]), .c_out(c[35]));
    fullAdder fa32 (.a(mode == 2'b01 ? 1'b1 : p[03][13]), .b(p[04][11]), .c_in(p[05][09]), .s(s[36]), .c_out(c[36]));
    fullAdder fa33 (.a(p[06][07]), .b(p[07][05]), .c_in(p[08][03]), .s(s[37]), .c_out(c[37]));
    fullAdder fa34 (.a(p[00][20]), .b(p[01][18]), .c_in(p[02][16]), .s(s[38]), .c_out(c[38]));
    fullAdder fa35 (.a(p[03][14]), .b(mode == 2'b01 ? ~comp[4] : p[04][12]), .c_in(p[05][10]), .s(s[39]), .c_out(c[39]));
    fullAdder fa36 (.a(p[06][08]), .b(p[07][06]), .c_in(p[08][04]), .s(s[40]), .c_out(c[40]));
    fullAdder fa37 (.a(p[09][02]), .b(p[10][00]), .c_in(mode == 2'b01 ? 1'b0 : comp[10]), .s(s[41]), .c_out(c[41]));
    fullAdder fa38 (.a(p[00][21]), .b(p[01][19]), .c_in(p[02][17]), .s(s[42]), .c_out(c[42]));
    fullAdder fa39 (.a(p[03][15]), .b(mode == 2'b01 ? 1'b1 : p[04][13]), .c_in(p[05][11]), .s(s[43]), .c_out(c[43]));
    fullAdder fa40 (.a(p[06][09]), .b(p[07][07]), .c_in(p[08][05]), .s(s[44]), .c_out(c[44]));
    halfAdder ha6 (.a(p[09][03]), .b(p[10][01]), .s(s[45]), .c_out(c[45]));
    fullAdder fa41 (.a(p[00][22]), .b(p[01][20]), .c_in(p[02][18]), .s(s[46]), .c_out(c[46]));
    fullAdder fa42 (.a(p[03][16]), .b(p[04][14]), .c_in(p[05][12]), .s(s[47]), .c_out(c[47]));
    fullAdder fa43 (.a(p[06][10]), .b(p[07][08]), .c_in(p[08][06]), .s(s[48]), .c_out(c[48]));
    fullAdder fa44 (.a(p[09][04]), .b(p[10][02]), .c_in(p[11][00]), .s(s[49]), .c_out(c[49]));
    fullAdder fa45 (.a(p[00][23]), .b(p[01][21]), .c_in(p[02][19]), .s(s[50]), .c_out(c[50]));
    fullAdder fa46 (.a(p[03][17]), .b(p[04][15]), .c_in(p[05][13]), .s(s[51]), .c_out(c[51]));
    fullAdder fa47 (.a(p[06][11]), .b(p[07][09]), .c_in(p[08][07]), .s(s[52]), .c_out(c[52]));
    fullAdder fa48 (.a(p[09][05]), .b(p[10][03]), .c_in(p[11][01]), .s(s[53]), .c_out(c[53]));
    fullAdder fa49 (.a(p[00][24]), .b(p[01][22]), .c_in(p[02][20]), .s(s[54]), .c_out(c[54]));
    fullAdder fa50 (.a(p[03][18]), .b(p[04][16]), .c_in(p[05][14]), .s(s[55]), .c_out(c[55]));
    fullAdder fa51 (.a(p[06][12]), .b(p[07][10]), .c_in(p[08][08]), .s(s[56]), .c_out(c[56]));
    fullAdder fa52 (.a(p[09][06]), .b(p[10][04]), .c_in(p[11][02]), .s(s[57]), .c_out(c[57]));
    halfAdder ha7 (.a(p[12][00]), .b(mode == 2'b11 ?  comp[12] : 1'b0), .s(s[58]), .c_out(c[58]));
    fullAdder fa53 (.a(mode == 2'b10 ? comp[0] : p[00][25]), .b(p[01][23]), .c_in(p[02][21]), .s(s[59]), .c_out(c[59]));
    fullAdder fa54 (.a(p[03][19]), .b(p[04][17]), .c_in(p[05][15]), .s(s[60]), .c_out(c[60]));
    fullAdder fa55 (.a(p[06][13]), .b(p[07][11]), .c_in(p[08][09]), .s(s[61]), .c_out(c[61]));
    fullAdder fa56 (.a(p[09][07]), .b(p[10][05]), .c_in(p[11][03]), .s(s[62]), .c_out(c[62]));
    fullAdder fa57 (.a(mode == 2'b10 ? comp[0] : p[00][26]), .b(p[01][24]), .c_in(p[02][22]), .s(s[63]), .c_out(c[63]));
    fullAdder fa58 (.a(p[03][20]), .b(p[04][18]), .c_in(p[05][16]), .s(s[64]), .c_out(c[64]));
    fullAdder fa59 (.a(p[06][14]), .b(p[07][12]), .c_in(p[08][10]), .s(s[65]), .c_out(c[65]));
    fullAdder fa60 (.a(p[09][08]), .b(p[10][06]), .c_in(p[11][04]), .s(s[66]), .c_out(c[66]));
    fullAdder fa61 (.a(p[12][02]), .b(p[13][00]), .c_in(mode == 2'b11 ?  comp[13] : 1'b0), .s(s[67]), .c_out(c[67]));
    fullAdder fa62 (.a(mode == 2'b10 ? ~comp[0] : p[00][27]), .b(mode == 2'b10 ? ~comp[1] : p[01][25]), .c_in(p[02][23]), .s(s[68]), .c_out(c[68]));
    fullAdder fa63 (.a(p[03][21]), .b(p[04][19]), .c_in(p[05][17]), .s(s[69]), .c_out(c[69]));
    fullAdder fa64 (.a(p[06][15]), .b(p[07][13]), .c_in(p[08][11]), .s(s[70]), .c_out(c[70]));
    fullAdder fa65 (.a(p[09][09]), .b(p[10][07]), .c_in(p[11][05]), .s(s[71]), .c_out(c[71]));
    halfAdder ha8 (.a(p[12][03]), .b(p[13][01]), .s(s[72]), .c_out(c[72]));
    fullAdder fa66 (.a(p[00][28]), .b(mode == 2'b10 ? 1'b1 : p[01][26]), .c_in(p[02][24]), .s(s[73]), .c_out(c[73]));
    fullAdder fa67 (.a(p[03][22]), .b(p[04][20]), .c_in(p[05][18]), .s(s[74]), .c_out(c[74]));
    fullAdder fa68 (.a(p[06][16]), .b(p[07][14]), .c_in(mode == 2'b01 ? comp[7] : p[08][12]), .s(s[75]), .c_out(c[75]));
    fullAdder fa69 (.a(p[09][10]), .b(p[10][08]), .c_in(p[11][06]), .s(s[76]), .c_out(c[76]));
    fullAdder fa70 (.a(p[12][04]), .b(p[13][02]), .c_in(p[14][00]), .s(s[77]), .c_out(c[77]));
    fullAdder fa71 (.a(p[00][29]), .b(p[01][27]), .c_in(mode == 2'b10 ? ~comp[2] : p[02][25]), .s(s[78]), .c_out(c[78]));
    fullAdder fa72 (.a(p[03][23]), .b(p[04][21]), .c_in(p[05][19]), .s(s[79]), .c_out(c[79]));
    fullAdder fa73 (.a(p[06][17]), .b(p[07][15]), .c_in(p[08][13]), .s(s[80]), .c_out(c[80]));
    fullAdder fa74 (.a(p[09][11]), .b(p[10][09]), .c_in(p[11][07]), .s(s[81]), .c_out(c[81]));
    fullAdder fa75 (.a(p[12][05]), .b(p[13][03]), .c_in(p[14][01]), .s(s[82]), .c_out(c[82]));
    fullAdder fa76 (.a(p[00][30]), .b(p[01][28]), .c_in(mode == 2'b10 ? 1'b1 : p[02][26]), .s(s[83]), .c_out(c[83]));
    fullAdder fa77 (.a(p[03][24]), .b(p[04][22]), .c_in(p[05][20]), .s(s[84]), .c_out(c[84]));
    fullAdder fa78 (.a(p[06][18]), .b(p[07][16]), .c_in(p[08][14]), .s(s[85]), .c_out(c[85]));
    fullAdder fa79 (.a(mode == 2'b01 ? comp[8] : p[09][12]), .b(p[10][10]), .c_in(p[11][08]), .s(s[86]), .c_out(c[86]));
    fullAdder fa80 (.a(p[12][06]), .b(p[13][04]), .c_in(p[14][02]), .s(s[87]), .c_out(c[87]));
    halfAdder ha9 (.a(p[15][00]), .b(mode == 2'b11 ? comp[15] : 1'b0), .s(s[88]), .c_out(c[88]));
    fullAdder fa81 (.a(p[00][31]), .b(p[01][29]), .c_in(p[02][27]), .s(s[89]), .c_out(c[89]));
    fullAdder fa82 (.a(mode == 2'b10 ? ~comp[3] : p[03][25]), .b(p[04][23]), .c_in(p[05][21]), .s(s[90]), .c_out(c[90]));
    fullAdder fa83 (.a(p[06][19]), .b(p[07][17]), .c_in(p[08][15]), .s(s[91]), .c_out(c[91]));
    fullAdder fa84 (.a(p[09][13]), .b(p[10][11]), .c_in(p[11][09]), .s(s[92]), .c_out(c[92]));
    fullAdder fa85 (.a(p[12][07]), .b(p[13][05]), .c_in(p[14][03]), .s(s[93]), .c_out(c[93]));
    fullAdder fa86 (.a(p[00][32]), .b(p[01][30]), .c_in(p[02][28]), .s(s[94]), .c_out(c[94]));
    fullAdder fa87 (.a(mode == 2'b10 ? 1'b1 : p[03][26]), .b(p[04][24]), .c_in(p[05][22]), .s(s[95]), .c_out(c[95]));
    fullAdder fa88 (.a(p[06][20]), .b(p[07][18]), .c_in(p[08][16]), .s(s[96]), .c_out(c[96]));
    fullAdder fa89 (.a(p[09][14]), .b(mode == 2'b01 ? comp[9] : p[10][12]), .c_in(p[11][10]), .s(s[97]), .c_out(c[97]));
    fullAdder fa90 (.a(p[12][08]), .b(p[13][06]), .c_in(p[14][04]), .s(s[98]), .c_out(c[98]));
    fullAdder fa91 (.a(p[15][02]), .b(p[16][00]), .c_in(mode == 2'b11 ? comp[16] : 1'b0), .s(s[99]), .c_out(c[99]));
    fullAdder fa92 (.a(p[00][33]), .b(p[01][31]), .c_in(p[02][29]), .s(s[100]), .c_out(c[100]));
    fullAdder fa93 (.a(p[03][27]), .b(mode == 2'b10 ? ~comp[4] : p[04][25]), .c_in(p[05][23]), .s(s[101]), .c_out(c[101]));
    fullAdder fa94 (.a(p[06][21]), .b(p[07][19]), .c_in(p[08][17]), .s(s[102]), .c_out(c[102]));
    fullAdder fa95 (.a(p[09][15]), .b(p[10][13]), .c_in(p[11][11]), .s(s[103]), .c_out(c[103]));
    fullAdder fa96 (.a(p[12][09]), .b(p[13][07]), .c_in(p[14][05]), .s(s[104]), .c_out(c[104]));
    halfAdder ha10 (.a(p[15][03]), .b(p[16][01]), .s(s[105]), .c_out(c[105]));
    fullAdder fa97 (.a(p[00][34]), .b(p[01][32]), .c_in(p[02][30]), .s(s[106]), .c_out(c[106]));
    fullAdder fa98 (.a(p[03][28]), .b(mode == 2'b10 ? 1'b1 : p[04][26]), .c_in(p[05][24]), .s(s[107]), .c_out(c[107]));
    fullAdder fa99 (.a(p[06][22]), .b(p[07][20]), .c_in(p[08][18]), .s(s[108]), .c_out(c[108]));
    fullAdder fa100 (.a(p[09][16]), .b(p[10][14]), .c_in(mode == 2'b01 ? comp[10] : p[11][12]), .s(s[109]), .c_out(c[109]));
    fullAdder fa101 (.a(p[12][10]), .b(p[13][08]), .c_in(p[14][06]), .s(s[110]), .c_out(c[110]));
    fullAdder fa102 (.a(p[15][04]), .b(p[16][02]), .c_in(p[17][00]), .s(s[111]), .c_out(c[111]));
    fullAdder fa103 (.a(p[00][35]), .b(p[01][33]), .c_in(p[02][31]), .s(s[112]), .c_out(c[112]));
    fullAdder fa104 (.a(p[03][29]), .b(p[04][27]), .c_in(mode == 2'b10 ? ~comp[5] : p[05][25]), .s(s[113]), .c_out(c[113]));
    fullAdder fa105 (.a(p[06][23]), .b(p[07][21]), .c_in(p[08][19]), .s(s[114]), .c_out(c[114]));
    fullAdder fa106 (.a(p[09][17]), .b(p[10][15]), .c_in(p[11][13]), .s(s[115]), .c_out(c[115]));
    fullAdder fa107 (.a(p[12][11]), .b(p[13][09]), .c_in(p[14][07]), .s(s[116]), .c_out(c[116]));
    fullAdder fa108 (.a(p[15][05]), .b(p[16][03]), .c_in(p[17][01]), .s(s[117]), .c_out(c[117]));
    fullAdder fa109 (.a(p[00][36]), .b(p[01][34]), .c_in(p[02][32]), .s(s[118]), .c_out(c[118]));
    fullAdder fa110 (.a(p[03][30]), .b(p[04][28]), .c_in(mode == 2'b10 ? 1'b1 : p[05][26]), .s(s[119]), .c_out(c[119]));
    fullAdder fa111 (.a(p[06][24]), .b(p[07][22]), .c_in(p[08][20]), .s(s[120]), .c_out(c[120]));
    fullAdder fa112 (.a(p[09][18]), .b(p[10][16]), .c_in(p[11][14]), .s(s[121]), .c_out(c[121]));
    fullAdder fa113 (.a(mode == 2'b01 ? comp[11] : p[12][12]), .b(p[13][10]), .c_in(p[14][08]), .s(s[122]), .c_out(c[122]));
    fullAdder fa114 (.a(p[15][06]), .b(p[16][04]), .c_in(p[17][02]), .s(s[123]), .c_out(c[123]));
    halfAdder ha11 (.a(p[18][00]), .b(mode == 2'b11 ? comp[18] : 1'b0), .s(s[124]), .c_out(c[124]));
    fullAdder fa115 (.a(p[00][37]), .b(p[01][35]), .c_in(p[02][33]), .s(s[125]), .c_out(c[125]));
    fullAdder fa116 (.a(p[03][31]), .b(p[04][29]), .c_in(p[05][27]), .s(s[126]), .c_out(c[126]));
    fullAdder fa117 (.a(mode == 2'b10 ? ~comp[6] : p[06][25]), .b(p[07][23]), .c_in(p[08][21]), .s(s[127]), .c_out(c[127]));
    fullAdder fa118 (.a(p[09][19]), .b(p[10][17]), .c_in(p[11][15]), .s(s[128]), .c_out(c[128]));
    fullAdder fa119 (.a(p[12][13]), .b(p[13][11]), .c_in(p[14][09]), .s(s[129]), .c_out(c[129]));
    fullAdder fa120 (.a(p[15][07]), .b(p[16][05]), .c_in(p[17][03]), .s(s[130]), .c_out(c[130]));
    fullAdder fa121 (.a(p[00][38]), .b(p[01][36]), .c_in(p[02][34]), .s(s[131]), .c_out(c[131]));
    fullAdder fa122 (.a(p[03][32]), .b(p[04][30]), .c_in(p[05][28]), .s(s[132]), .c_out(c[132]));
    fullAdder fa123 (.a(mode == 2'b10 ? 1'b1 : p[06][26]), .b(p[07][24]), .c_in(p[08][22]), .s(s[133]), .c_out(c[133]));
    fullAdder fa124 (.a(p[09][20]), .b(p[10][18]), .c_in(p[11][16]), .s(s[134]), .c_out(c[134]));
    fullAdder fa125 (.a(p[12][14]), .b(p[13][12]), .c_in(p[14][10]), .s(s[135]), .c_out(c[135]));
    fullAdder fa126 (.a(p[15][08]), .b(p[16][06]), .c_in(p[17][04]), .s(s[136]), .c_out(c[136]));
    fullAdder fa127 (.a(p[18][02]), .b(p[19][00]), .c_in(mode == 2'b11 ? comp[19] : 1'b0), .s(s[137]), .c_out(c[137]));
    fullAdder fa128 (.a(p[00][39]), .b(p[01][37]), .c_in(p[02][35]), .s(s[138]), .c_out(c[138]));
    fullAdder fa129 (.a(p[03][33]), .b(p[04][31]), .c_in(p[05][29]), .s(s[139]), .c_out(c[139]));
    fullAdder fa130 (.a(p[06][27]), .b(mode == 2'b10 ? ~comp[7] : p[07][25]), .c_in(p[08][23]), .s(s[140]), .c_out(c[140]));
    fullAdder fa131 (.a(p[09][21]), .b(p[10][19]), .c_in(p[11][17]), .s(s[141]), .c_out(c[141]));
    fullAdder fa132 (.a(p[12][15]), .b(p[13][13]), .c_in(p[14][11]), .s(s[142]), .c_out(c[142]));
    fullAdder fa133 (.a(p[15][09]), .b(p[16][07]), .c_in(p[17][05]), .s(s[143]), .c_out(c[143]));
    halfAdder ha12 (.a(p[18][03]), .b(p[19][01]), .s(s[144]), .c_out(c[144]));
    fullAdder fa134 (.a(p[00][40]), .b(p[01][38]), .c_in(p[02][36]), .s(s[145]), .c_out(c[145]));
    fullAdder fa135 (.a(p[03][34]), .b(p[04][32]), .c_in(p[05][30]), .s(s[146]), .c_out(c[146]));
    fullAdder fa136 (.a(p[06][28]), .b(mode == 2'b10 ? 1'b1 : mode == 2'b01 ? comp[7] : p[07][26]), .c_in(p[08][24]), .s(s[147]), .c_out(c[147]));
    fullAdder fa137 (.a(p[09][22]), .b(p[10][20]), .c_in(p[11][18]), .s(s[148]), .c_out(c[148]));
    fullAdder fa138 (.a(p[12][16]), .b(p[13][14]), .c_in(p[14][12]), .s(s[149]), .c_out(c[149]));
    fullAdder fa139 (.a(p[15][10]), .b(p[16][08]), .c_in(p[17][06]), .s(s[150]), .c_out(c[150]));
    fullAdder fa140 (.a(p[18][04]), .b(p[19][02]), .c_in(p[20][00]), .s(s[151]), .c_out(c[151]));
    fullAdder fa141 (.a(p[00][41]), .b(p[01][39]), .c_in(p[02][37]), .s(s[152]), .c_out(c[152]));
    fullAdder fa142 (.a(p[03][35]), .b(p[04][33]), .c_in(p[05][31]), .s(s[153]), .c_out(c[153]));
    fullAdder fa143 (.a(p[06][29]), .b(mode == 2'b01 ? comp[7] : p[07][27]), .c_in(mode == 2'b10 ? ~comp[8] : p[08][25]), .s(s[154]), .c_out(c[154]));
    fullAdder fa144 (.a(p[09][23]), .b(p[10][21]), .c_in(p[11][19]), .s(s[155]), .c_out(c[155]));
    fullAdder fa145 (.a(p[12][17]), .b(p[13][15]), .c_in(p[14][13]), .s(s[156]), .c_out(c[156]));
    fullAdder fa146 (.a(p[15][11]), .b(p[16][09]), .c_in(p[17][07]), .s(s[157]), .c_out(c[157]));
    fullAdder fa147 (.a(p[18][05]), .b(p[19][03]), .c_in(p[20][01]), .s(s[158]), .c_out(c[158]));
    fullAdder fa148 (.a(p[00][42]), .b(p[01][40]), .c_in(p[02][38]), .s(s[159]), .c_out(c[159]));
    fullAdder fa149 (.a(p[03][36]), .b(p[04][34]), .c_in(p[05][32]), .s(s[160]), .c_out(c[160]));
    fullAdder fa150 (.a(p[06][30]), .b(mode == 2'b01 ? ~comp[7] : p[07][28]), .c_in(mode == 2'b10 ? 1'b1 : mode == 2'b01 ? ~comp[8] : p[08][26]), .s(s[161]), .c_out(c[161]));
    fullAdder fa151 (.a(p[09][24]), .b(p[10][22]), .c_in(p[11][20]), .s(s[162]), .c_out(c[162]));
    fullAdder fa152 (.a(p[12][18]), .b(p[13][16]), .c_in(p[14][14]), .s(s[163]), .c_out(c[163]));
    fullAdder fa153 (.a(p[15][12]), .b(p[16][10]), .c_in(p[17][08]), .s(s[164]), .c_out(c[164]));
    fullAdder fa154 (.a(p[18][06]), .b(p[19][04]), .c_in(p[20][02]), .s(s[165]), .c_out(c[165]));
    halfAdder ha13 (.a(p[21][00]), .b(mode == 2'b11 ? comp[21] : 1'b0), .s(s[166]), .c_out(c[166]));
    fullAdder fa155 (.a(p[00][43]), .b(p[01][41]), .c_in(p[02][39]), .s(s[167]), .c_out(c[167]));
    fullAdder fa156 (.a(p[03][37]), .b(p[04][35]), .c_in(p[05][33]), .s(s[168]), .c_out(c[168]));
    fullAdder fa157 (.a(p[06][31]), .b(p[07][29]), .c_in(mode == 2'b01 ? 1'b1 : p[08][27]), .s(s[169]), .c_out(c[169]));
    fullAdder fa158 (.a(mode == 2'b10 ? ~comp[9] : p[09][25]), .b(p[10][23]), .c_in(p[11][21]), .s(s[170]), .c_out(c[170]));
    fullAdder fa159 (.a(p[12][19]), .b(p[13][17]), .c_in(p[14][15]), .s(s[171]), .c_out(c[171]));
    fullAdder fa160 (.a(p[15][13]), .b(p[16][11]), .c_in(p[17][09]), .s(s[172]), .c_out(c[172]));
    fullAdder fa161 (.a(p[18][07]), .b(p[19][05]), .c_in(p[20][03]), .s(s[173]), .c_out(c[173]));
    fullAdder fa162 (.a(p[00][44]), .b(p[01][42]), .c_in(p[02][40]), .s(s[174]), .c_out(c[174]));
    fullAdder fa163 (.a(p[03][38]), .b(p[04][36]), .c_in(p[05][34]), .s(s[175]), .c_out(c[175]));
    fullAdder fa164 (.a(p[06][32]), .b(p[07][30]), .c_in(p[08][28]), .s(s[176]), .c_out(c[176]));
    fullAdder fa165 (.a(mode == 2'b10 ? 1'b1 : mode == 2'b01 ? ~comp[9] : p[09][26]), .b(p[10][24]), .c_in(p[11][22]), .s(s[177]), .c_out(c[177]));
    fullAdder fa166 (.a(p[12][20]), .b(p[13][18]), .c_in(p[14][16]), .s(s[178]), .c_out(c[178]));
    fullAdder fa167 (.a(p[15][14]), .b(p[16][12]), .c_in(p[17][10]), .s(s[179]), .c_out(c[179]));
    fullAdder fa168 (.a(p[18][08]), .b(p[19][06]), .c_in(p[20][04]), .s(s[180]), .c_out(c[180]));
    fullAdder fa169 (.a(p[21][02]), .b(p[22][00]), .c_in(mode == 2'b11 ? comp[22] : 1'b0), .s(s[181]), .c_out(c[181]));
    fullAdder fa170 (.a(p[00][45]), .b(p[01][43]), .c_in(p[02][41]), .s(s[182]), .c_out(c[182]));
    fullAdder fa171 (.a(p[03][39]), .b(p[04][37]), .c_in(p[05][35]), .s(s[183]), .c_out(c[183]));
    fullAdder fa172 (.a(p[06][33]), .b(p[07][31]), .c_in(p[08][29]), .s(s[184]), .c_out(c[184]));
    fullAdder fa173 (.a(mode == 2'b01 ? 1'b1 : p[09][27]), .b(mode == 2'b10 ? ~comp[10] : p[10][25]), .c_in(p[11][23]), .s(s[185]), .c_out(c[185]));
    fullAdder fa174 (.a(p[12][21]), .b(p[13][19]), .c_in(p[14][17]), .s(s[186]), .c_out(c[186]));
    fullAdder fa175 (.a(p[15][15]), .b(p[16][13]), .c_in(p[17][11]), .s(s[187]), .c_out(c[187]));
    fullAdder fa176 (.a(p[18][09]), .b(p[19][07]), .c_in(p[20][05]), .s(s[188]), .c_out(c[188]));
    halfAdder ha14 (.a(p[21][03]), .b(p[22][01]), .s(s[189]), .c_out(c[189]));
    fullAdder fa177 (.a(p[00][46]), .b(p[01][44]), .c_in(p[02][42]), .s(s[190]), .c_out(c[190]));
    fullAdder fa178 (.a(p[03][40]), .b(p[04][38]), .c_in(p[05][36]), .s(s[191]), .c_out(c[191]));
    fullAdder fa179 (.a(p[06][34]), .b(p[07][32]), .c_in(p[08][30]), .s(s[192]), .c_out(c[192]));
    fullAdder fa180 (.a(p[09][28]), .b(mode == 2'b10 ? 1'b1 : mode == 2'b01 ? ~comp[10] : p[10][26]), .c_in(p[11][24]), .s(s[193]), .c_out(c[193]));
    fullAdder fa181 (.a(p[12][22]), .b(p[13][20]), .c_in(p[14][18]), .s(s[194]), .c_out(c[194]));
    fullAdder fa182 (.a(p[15][16]), .b(p[16][14]), .c_in(p[17][12]), .s(s[195]), .c_out(c[195]));
    fullAdder fa183 (.a(p[18][10]), .b(p[19][08]), .c_in(p[20][06]), .s(s[196]), .c_out(c[196]));
    fullAdder fa184 (.a(p[21][04]), .b(p[22][02]), .c_in(p[23][00]), .s(s[197]), .c_out(c[197]));
    fullAdder fa185 (.a(p[00][47]), .b(p[01][45]), .c_in(p[02][43]), .s(s[198]), .c_out(c[198]));
    fullAdder fa186 (.a(p[03][41]), .b(p[04][39]), .c_in(p[05][37]), .s(s[199]), .c_out(c[199]));
    fullAdder fa187 (.a(p[06][35]), .b(p[07][33]), .c_in(p[08][31]), .s(s[200]), .c_out(c[200]));
    fullAdder fa188 (.a(p[09][29]), .b(mode == 2'b01 ? 1'b1 : p[10][27]), .c_in(mode == 2'b10 ? ~comp[11] : p[11][25]), .s(s[201]), .c_out(c[201]));
    fullAdder fa189 (.a(p[12][23]), .b(p[13][21]), .c_in(p[14][19]), .s(s[202]), .c_out(c[202]));
    fullAdder fa190 (.a(p[15][17]), .b(p[16][15]), .c_in(p[17][13]), .s(s[203]), .c_out(c[203]));
    fullAdder fa191 (.a(p[18][11]), .b(p[19][09]), .c_in(p[20][07]), .s(s[204]), .c_out(c[204]));
    fullAdder fa192 (.a(p[21][05]), .b(p[22][03]), .c_in(p[23][01]), .s(s[205]), .c_out(c[205]));
    fullAdder fa193 (.a(p[00][48]), .b(p[01][46]), .c_in(p[02][44]), .s(s[206]), .c_out(c[206]));
    fullAdder fa194 (.a(p[03][42]), .b(p[04][40]), .c_in(p[05][38]), .s(s[207]), .c_out(c[207]));
    fullAdder fa195 (.a(p[06][36]), .b(p[07][34]), .c_in(p[08][32]), .s(s[208]), .c_out(c[208]));
    fullAdder fa196 (.a(p[09][30]), .b(p[10][28]), .c_in(mode == 2'b01 ? ~comp[11] : p[11][26]), .s(s[209]), .c_out(c[209]));
    fullAdder fa197 (.a(mode == 2'b10 ? 1'b0 : p[12][24]), .b(p[13][22]), .c_in(p[14][20]), .s(s[210]), .c_out(c[210]));
    fullAdder fa198 (.a(p[15][18]), .b(p[16][16]), .c_in(p[17][14]), .s(s[211]), .c_out(c[211]));
    fullAdder fa199 (.a(p[18][12]), .b(p[19][10]), .c_in(p[20][08]), .s(s[212]), .c_out(c[212]));
    fullAdder fa200 (.a(p[21][06]), .b(p[22][04]), .c_in(p[23][02]), .s(s[213]), .c_out(c[213]));
    halfAdder ha15 (.a(p[24][00]), .b(mode == 2'b11 ? comp[24] : 1'b0), .s(s[214]), .c_out(c[214]));
    fullAdder fa201 (.a(p[00][49]), .b(p[01][47]), .c_in(p[02][45]), .s(s[215]), .c_out(c[215]));
    fullAdder fa202 (.a(p[03][43]), .b(p[04][41]), .c_in(p[05][39]), .s(s[216]), .c_out(c[216]));
    fullAdder fa203 (.a(p[06][37]), .b(p[07][35]), .c_in(p[08][33]), .s(s[217]), .c_out(c[217]));
    fullAdder fa204 (.a(p[09][31]), .b(p[10][29]), .c_in(mode == 2'b01 ? 1'b1 : p[11][27]), .s(s[218]), .c_out(c[218]));
    fullAdder fa205 (.a(p[12][25]), .b(p[13][23]), .c_in(p[14][21]), .s(s[219]), .c_out(c[219]));
    fullAdder fa206 (.a(p[15][19]), .b(p[16][17]), .c_in(p[17][15]), .s(s[220]), .c_out(c[220]));
    fullAdder fa207 (.a(p[18][13]), .b(p[19][11]), .c_in(p[20][09]), .s(s[221]), .c_out(c[221]));
    fullAdder fa208 (.a(p[21][07]), .b(p[22][05]), .c_in(p[23][03]), .s(s[222]), .c_out(c[222]));
    fullAdder fa209 (.a(p[00][50]), .b(p[01][48]), .c_in(p[02][46]), .s(s[223]), .c_out(c[223]));
    fullAdder fa210 (.a(p[03][44]), .b(p[04][42]), .c_in(p[05][40]), .s(s[224]), .c_out(c[224]));
    fullAdder fa211 (.a(p[06][38]), .b(p[07][36]), .c_in(p[08][34]), .s(s[225]), .c_out(c[225]));
    fullAdder fa212 (.a(p[09][32]), .b(p[10][30]), .c_in(p[11][28]), .s(s[226]), .c_out(c[226]));
    fullAdder fa213 (.a(p[12][26]), .b(p[13][24]), .c_in(p[14][22]), .s(s[227]), .c_out(c[227]));
    fullAdder fa214 (.a(p[15][20]), .b(p[16][18]), .c_in(p[17][16]), .s(s[228]), .c_out(c[228]));
    fullAdder fa215 (.a(p[18][14]), .b(p[19][12]), .c_in(p[20][10]), .s(s[229]), .c_out(c[229]));
    fullAdder fa216 (.a(p[21][08]), .b(p[22][06]), .c_in(p[23][04]), .s(s[230]), .c_out(c[230]));
    fullAdder fa217 (.a(p[24][02]), .b(p[25][00]), .c_in(mode == 2'b11 ? comp[25] : 1'b0), .s(s[231]), .c_out(c[231]));
    fullAdder fa218 (.a(p[00][51]), .b(p[01][49]), .c_in(p[02][47]), .s(s[232]), .c_out(c[232]));
    fullAdder fa219 (.a(p[03][45]), .b(p[04][43]), .c_in(p[05][41]), .s(s[233]), .c_out(c[233]));
    fullAdder fa220 (.a(p[06][39]), .b(p[07][37]), .c_in(p[08][35]), .s(s[234]), .c_out(c[234]));
    fullAdder fa221 (.a(p[09][33]), .b(p[10][31]), .c_in(p[11][29]), .s(s[235]), .c_out(c[235]));
    fullAdder fa222 (.a(p[12][27]), .b(p[13][25]), .c_in(p[14][23]), .s(s[236]), .c_out(c[236]));
    fullAdder fa223 (.a(p[15][21]), .b(p[16][19]), .c_in(p[17][17]), .s(s[237]), .c_out(c[237]));
    fullAdder fa224 (.a(p[18][15]), .b(p[19][13]), .c_in(p[20][11]), .s(s[238]), .c_out(c[238]));
    fullAdder fa225 (.a(p[21][09]), .b(p[22][07]), .c_in(p[23][05]), .s(s[239]), .c_out(c[239]));
    halfAdder ha16 (.a(p[24][03]), .b(p[25][01]), .s(s[240]), .c_out(c[240]));
    fullAdder fa226 (.a(p[00][52]), .b(p[01][50]), .c_in(p[02][48]), .s(s[241]), .c_out(c[241]));
    fullAdder fa227 (.a(p[03][46]), .b(p[04][44]), .c_in(p[05][42]), .s(s[242]), .c_out(c[242]));
    fullAdder fa228 (.a(p[06][40]), .b(p[07][38]), .c_in(p[08][36]), .s(s[243]), .c_out(c[243]));
    fullAdder fa229 (.a(p[09][34]), .b(p[10][32]), .c_in(p[11][30]), .s(s[244]), .c_out(c[244]));
    fullAdder fa230 (.a(p[12][28]), .b(p[13][26]), .c_in(p[14][24]), .s(s[245]), .c_out(c[245]));
    fullAdder fa231 (.a(p[15][22]), .b(p[16][20]), .c_in(p[17][18]), .s(s[246]), .c_out(c[246]));
    fullAdder fa232 (.a(p[18][16]), .b(p[19][14]), .c_in(p[20][12]), .s(s[247]), .c_out(c[247]));
    fullAdder fa233 (.a(p[21][10]), .b(p[22][08]), .c_in(p[23][06]), .s(s[248]), .c_out(c[248]));
    fullAdder fa234 (.a(p[24][04]), .b(p[25][02]), .c_in(p[26][00]), .s(s[249]), .c_out(c[249]));
    fullAdder fa235 (.a(p[00][53]), .b(p[01][51]), .c_in(p[02][49]), .s(s[250]), .c_out(c[250]));
    fullAdder fa236 (.a(p[03][47]), .b(p[04][45]), .c_in(p[05][43]), .s(s[251]), .c_out(c[251]));
    fullAdder fa237 (.a(p[06][41]), .b(p[07][39]), .c_in(p[08][37]), .s(s[252]), .c_out(c[252]));
    fullAdder fa238 (.a(p[09][35]), .b(p[10][33]), .c_in(p[11][31]), .s(s[253]), .c_out(c[253]));
    fullAdder fa239 (.a(p[12][29]), .b(p[13][27]), .c_in(p[14][25]), .s(s[254]), .c_out(c[254]));
    fullAdder fa240 (.a(p[15][23]), .b(p[16][21]), .c_in(p[17][19]), .s(s[255]), .c_out(c[255]));
    fullAdder fa241 (.a(p[18][17]), .b(p[19][15]), .c_in(p[20][13]), .s(s[256]), .c_out(c[256]));
    fullAdder fa242 (.a(p[21][11]), .b(p[22][09]), .c_in(p[23][07]), .s(s[257]), .c_out(c[257]));
    fullAdder fa243 (.a(p[24][05]), .b(p[25][03]), .c_in(p[26][01]), .s(s[258]), .c_out(c[258]));
    fullAdder fa244 (.a(mode == 2'b11 ? comp[0] : 1'b0), .b(p[01][52]), .c_in(p[02][50]), .s(s[259]), .c_out(c[259]));
    fullAdder fa245 (.a(p[03][48]), .b(p[04][46]), .c_in(p[05][44]), .s(s[260]), .c_out(c[260]));
    fullAdder fa246 (.a(p[06][42]), .b(p[07][40]), .c_in(p[08][38]), .s(s[261]), .c_out(c[261]));
    fullAdder fa247 (.a(p[09][36]), .b(p[10][34]), .c_in(p[11][32]), .s(s[262]), .c_out(c[262]));
    fullAdder fa248 (.a(p[12][30]), .b(p[13][28]), .c_in(p[14][26]), .s(s[263]), .c_out(c[263]));
    fullAdder fa249 (.a(p[15][24]), .b(p[16][22]), .c_in(p[17][20]), .s(s[264]), .c_out(c[264]));
    fullAdder fa250 (.a(p[18][18]), .b(p[19][16]), .c_in(p[20][14]), .s(s[265]), .c_out(c[265]));
    fullAdder fa251 (.a(p[21][12]), .b(p[22][10]), .c_in(p[23][08]), .s(s[266]), .c_out(c[266]));
    fullAdder fa252 (.a(p[24][06]), .b(p[25][04]), .c_in(p[26][02]), .s(s[267]), .c_out(c[267]));
    fullAdder fa253 (.a(mode == 2'b11 ? comp[0] : 1'b0), .b(p[01][53]), .c_in(p[02][51]), .s(s[268]), .c_out(c[268]));
    fullAdder fa254 (.a(p[03][49]), .b(p[04][47]), .c_in(p[05][45]), .s(s[269]), .c_out(c[269]));
    fullAdder fa255 (.a(p[06][43]), .b(p[07][41]), .c_in(p[08][39]), .s(s[270]), .c_out(c[270]));
    fullAdder fa256 (.a(p[09][37]), .b(p[10][35]), .c_in(p[11][33]), .s(s[271]), .c_out(c[271]));
    fullAdder fa257 (.a(p[12][31]), .b(p[13][29]), .c_in(p[14][27]), .s(s[272]), .c_out(c[272]));
    fullAdder fa258 (.a(p[15][25]), .b(p[16][23]), .c_in(p[17][21]), .s(s[273]), .c_out(c[273]));
    fullAdder fa259 (.a(p[18][19]), .b(p[19][17]), .c_in(p[20][15]), .s(s[274]), .c_out(c[274]));
    fullAdder fa260 (.a(p[21][13]), .b(p[22][11]), .c_in(p[23][09]), .s(s[275]), .c_out(c[275]));
    fullAdder fa261 (.a(p[24][07]), .b(p[25][05]), .c_in(p[26][03]), .s(s[276]), .c_out(c[276]));
    fullAdder fa262 (.a(mode == 2'b11 ? ~comp[00] : 1'b0), .b(mode == 2'b11 ? ~comp[01] : 1'b0), .c_in(p[02][52]), .s(s[277]), .c_out(c[277]));
    fullAdder fa263 (.a(p[03][50]), .b(p[04][48]), .c_in(p[05][46]), .s(s[278]), .c_out(c[278]));
    fullAdder fa264 (.a(p[06][44]), .b(p[07][42]), .c_in(p[08][40]), .s(s[279]), .c_out(c[279]));
    fullAdder fa265 (.a(p[09][38]), .b(p[10][36]), .c_in(p[11][34]), .s(s[280]), .c_out(c[280]));
    fullAdder fa266 (.a(p[12][32]), .b(p[13][30]), .c_in(p[14][28]), .s(s[281]), .c_out(c[281]));
    fullAdder fa267 (.a(mode == 2'b01 ? comp[14] : p[15][26]), .b(p[16][24]), .c_in(p[17][22]), .s(s[282]), .c_out(c[282]));
    fullAdder fa268 (.a(p[18][20]), .b(p[19][18]), .c_in(p[20][16]), .s(s[283]), .c_out(c[283]));
    fullAdder fa269 (.a(p[21][14]), .b(p[22][12]), .c_in(p[23][10]), .s(s[284]), .c_out(c[284]));
    fullAdder fa270 (.a(p[24][08]), .b(p[25][06]), .c_in(p[26][04]), .s(s[285]), .c_out(c[285]));
    fullAdder fa271 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[02][53]), .c_in(p[03][51]), .s(s[286]), .c_out(c[286]));
    fullAdder fa272 (.a(p[04][49]), .b(p[05][47]), .c_in(p[06][45]), .s(s[287]), .c_out(c[287]));
    fullAdder fa273 (.a(p[07][43]), .b(p[08][41]), .c_in(p[09][39]), .s(s[288]), .c_out(c[288]));
    fullAdder fa274 (.a(p[10][37]), .b(p[11][35]), .c_in(p[12][33]), .s(s[289]), .c_out(c[289]));
    fullAdder fa275 (.a(p[13][31]), .b(p[14][29]), .c_in(mode == 2'b10 ? comp[14] : p[15][27]), .s(s[290]), .c_out(c[290]));
    fullAdder fa276 (.a(p[16][25]), .b(p[17][23]), .c_in(p[18][21]), .s(s[291]), .c_out(c[291]));
    fullAdder fa277 (.a(p[19][19]), .b(p[20][17]), .c_in(p[21][15]), .s(s[292]), .c_out(c[292]));
    fullAdder fa278 (.a(p[22][13]), .b(p[23][11]), .c_in(p[24][09]), .s(s[293]), .c_out(c[293]));
    halfAdder ha17 (.a(p[25][07]), .b(p[26][05]), .s(s[294]), .c_out(c[294]));
    fullAdder fa279 (.a(mode == 2'b11 ?  ~comp[02] : 1'b0), .b(p[03][52]), .c_in(p[04][50]), .s(s[295]), .c_out(c[295]));
    fullAdder fa280 (.a(p[05][48]), .b(p[06][46]), .c_in(p[07][44]), .s(s[296]), .c_out(c[296]));
    fullAdder fa281 (.a(p[08][42]), .b(p[09][40]), .c_in(p[10][38]), .s(s[297]), .c_out(c[297]));
    fullAdder fa282 (.a(p[11][36]), .b(p[12][34]), .c_in(p[13][32]), .s(s[298]), .c_out(c[298]));
    fullAdder fa283 (.a(p[14][30]), .b(p[15][28]), .c_in(mode == 2'b01 ? comp[15] : p[16][26]), .s(s[299]), .c_out(c[299]));
    fullAdder fa284 (.a(p[17][24]), .b(p[18][22]), .c_in(p[19][20]), .s(s[300]), .c_out(c[300]));
    fullAdder fa285 (.a(p[20][18]), .b(p[21][16]), .c_in(p[22][14]), .s(s[301]), .c_out(c[301]));
    fullAdder fa286 (.a(p[23][12]), .b(p[24][10]), .c_in(p[25][08]), .s(s[302]), .c_out(c[302]));
    fullAdder fa287 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[03][53]), .c_in(p[04][51]), .s(s[303]), .c_out(c[303]));
    fullAdder fa288 (.a(p[05][49]), .b(p[06][47]), .c_in(p[07][45]), .s(s[304]), .c_out(c[304]));
    fullAdder fa289 (.a(p[08][43]), .b(p[09][41]), .c_in(p[10][39]), .s(s[305]), .c_out(c[305]));
    fullAdder fa290 (.a(p[11][37]), .b(p[12][35]), .c_in(p[13][33]), .s(s[306]), .c_out(c[306]));
    fullAdder fa291 (.a(p[14][31]), .b(p[15][29]), .c_in(mode == 2'b10 ? comp[15] : p[16][27]), .s(s[307]), .c_out(c[307]));
    fullAdder fa292 (.a(p[17][25]), .b(p[18][23]), .c_in(p[19][21]), .s(s[308]), .c_out(c[308]));
    fullAdder fa293 (.a(p[20][19]), .b(p[21][17]), .c_in(p[22][15]), .s(s[309]), .c_out(c[309]));
    fullAdder fa294 (.a(p[23][13]), .b(p[24][11]), .c_in(p[25][09]), .s(s[310]), .c_out(c[310]));
    fullAdder fa295 (.a(mode == 2'b11 ?  ~comp[03] : 1'b0), .b(p[04][52]), .c_in(p[05][50]), .s(s[311]), .c_out(c[311]));
    fullAdder fa296 (.a(p[06][48]), .b(p[07][46]), .c_in(p[08][44]), .s(s[312]), .c_out(c[312]));
    fullAdder fa297 (.a(p[09][42]), .b(p[10][40]), .c_in(p[11][38]), .s(s[313]), .c_out(c[313]));
    fullAdder fa298 (.a(p[12][36]), .b(p[13][34]), .c_in(p[14][32]), .s(s[314]), .c_out(c[314]));
    fullAdder fa299 (.a(p[15][30]), .b(p[16][28]), .c_in(mode == 2'b01 ? comp[16] : p[17][26]), .s(s[315]), .c_out(c[315]));
    fullAdder fa300 (.a(p[18][24]), .b(p[19][22]), .c_in(p[20][20]), .s(s[316]), .c_out(c[316]));
    fullAdder fa301 (.a(p[21][18]), .b(p[22][16]), .c_in(p[23][14]), .s(s[317]), .c_out(c[317]));
    fullAdder fa302 (.a(p[24][12]), .b(p[25][10]), .c_in(p[26][08]), .s(s[318]), .c_out(c[318]));
    fullAdder fa303 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[04][53]), .c_in(p[05][51]), .s(s[319]), .c_out(c[319]));
    fullAdder fa304 (.a(p[06][49]), .b(p[07][47]), .c_in(p[08][45]), .s(s[320]), .c_out(c[320]));
    fullAdder fa305 (.a(p[09][43]), .b(p[10][41]), .c_in(p[11][39]), .s(s[321]), .c_out(c[321]));
    fullAdder fa306 (.a(p[12][37]), .b(p[13][35]), .c_in(p[14][33]), .s(s[322]), .c_out(c[322]));
    fullAdder fa307 (.a(p[15][31]), .b(p[16][29]), .c_in(mode == 2'b10 ? comp[16] : p[17][27]), .s(s[323]), .c_out(c[323]));
    fullAdder fa308 (.a(p[18][25]), .b(p[19][23]), .c_in(p[20][21]), .s(s[324]), .c_out(c[324]));
    fullAdder fa309 (.a(p[21][19]), .b(p[22][17]), .c_in(p[23][15]), .s(s[325]), .c_out(c[325]));
    fullAdder fa310 (.a(p[24][13]), .b(p[25][11]), .c_in(p[26][09]), .s(s[326]), .c_out(c[326]));
    fullAdder fa311 (.a(mode == 2'b11 ?  ~comp[04] : 1'b0), .b(p[05][52]), .c_in(p[06][50]), .s(s[327]), .c_out(c[327]));
    fullAdder fa312 (.a(p[07][48]), .b(p[08][46]), .c_in(p[09][44]), .s(s[328]), .c_out(c[328]));
    fullAdder fa313 (.a(p[10][42]), .b(p[11][40]), .c_in(p[12][38]), .s(s[329]), .c_out(c[329]));
    fullAdder fa314 (.a(p[13][36]), .b(p[14][34]), .c_in(p[15][32]), .s(s[330]), .c_out(c[330]));
    fullAdder fa315 (.a(p[16][30]), .b(p[17][28]), .c_in(mode == 2'b01 ? comp[17] : p[18][26]), .s(s[331]), .c_out(c[331]));
    fullAdder fa316 (.a(p[19][24]), .b(p[20][22]), .c_in(p[21][20]), .s(s[332]), .c_out(c[332]));
    fullAdder fa317 (.a(p[22][18]), .b(p[23][16]), .c_in(p[24][14]), .s(s[333]), .c_out(c[333]));
    halfAdder ha18 (.a(p[25][12]), .b(p[26][10]), .s(s[334]), .c_out(c[334]));
    fullAdder fa318 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[05][53]), .c_in(p[06][51]), .s(s[335]), .c_out(c[335]));
    fullAdder fa319 (.a(p[07][49]), .b(p[08][47]), .c_in(p[09][45]), .s(s[336]), .c_out(c[336]));
    fullAdder fa320 (.a(p[10][43]), .b(p[11][41]), .c_in(p[12][39]), .s(s[337]), .c_out(c[337]));
    fullAdder fa321 (.a(p[13][37]), .b(p[14][35]), .c_in(p[15][33]), .s(s[338]), .c_out(c[338]));
    fullAdder fa322 (.a(p[16][31]), .b(p[17][29]), .c_in(mode == 2'b10 ? comp[17] : p[18][27]), .s(s[339]), .c_out(c[339]));
    fullAdder fa323 (.a(p[19][25]), .b(p[20][23]), .c_in(p[21][21]), .s(s[340]), .c_out(c[340]));
    fullAdder fa324 (.a(p[22][19]), .b(p[23][17]), .c_in(p[24][15]), .s(s[341]), .c_out(c[341]));
    halfAdder ha19 (.a(p[25][13]), .b(p[26][11]), .s(s[342]), .c_out(c[342]));
    fullAdder fa325 (.a(mode == 2'b11 ?  ~comp[05] : 1'b0), .b(p[06][52]), .c_in(p[07][50]), .s(s[343]), .c_out(c[343]));
    fullAdder fa326 (.a(p[08][48]), .b(p[09][46]), .c_in(p[10][44]), .s(s[344]), .c_out(c[344]));
    fullAdder fa327 (.a(p[11][42]), .b(p[12][40]), .c_in(p[13][38]), .s(s[345]), .c_out(c[345]));
    fullAdder fa328 (.a(p[14][36]), .b(p[15][34]), .c_in(p[16][32]), .s(s[346]), .c_out(c[346]));
    fullAdder fa329 (.a(p[17][30]), .b(p[18][28]), .c_in(mode == 2'b01 ? comp[18] : p[19][26]), .s(s[347]), .c_out(c[347]));
    fullAdder fa330 (.a(p[20][24]), .b(p[21][22]), .c_in(p[22][20]), .s(s[348]), .c_out(c[348]));
    fullAdder fa331 (.a(p[23][18]), .b(p[24][16]), .c_in(p[25][14]), .s(s[349]), .c_out(c[349]));
    fullAdder fa332 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[06][53]), .c_in(p[07][51]), .s(s[350]), .c_out(c[350]));
    fullAdder fa333 (.a(p[08][49]), .b(p[09][47]), .c_in(p[10][45]), .s(s[351]), .c_out(c[351]));
    fullAdder fa334 (.a(p[11][43]), .b(p[12][41]), .c_in(p[13][39]), .s(s[352]), .c_out(c[352]));
    fullAdder fa335 (.a(p[14][37]), .b(p[15][35]), .c_in(p[16][33]), .s(s[353]), .c_out(c[353]));
    fullAdder fa336 (.a(p[17][31]), .b(p[18][29]), .c_in(mode == 2'b10 ? comp[18] : p[19][27]), .s(s[354]), .c_out(c[354]));
    fullAdder fa337 (.a(p[20][25]), .b(p[21][23]), .c_in(p[22][21]), .s(s[355]), .c_out(c[355]));
    fullAdder fa338 (.a(p[23][19]), .b(p[24][17]), .c_in(p[25][15]), .s(s[356]), .c_out(c[356]));
    fullAdder fa339 (.a(mode == 2'b11 ?  ~comp[06] : 1'b0), .b(p[07][52]), .c_in(p[08][50]), .s(s[357]), .c_out(c[357]));
    fullAdder fa340 (.a(p[09][48]), .b(p[10][46]), .c_in(p[11][44]), .s(s[358]), .c_out(c[358]));
    fullAdder fa341 (.a(p[12][42]), .b(p[13][40]), .c_in(p[14][38]), .s(s[359]), .c_out(c[359]));
    fullAdder fa342 (.a(p[15][36]), .b(p[16][34]), .c_in(p[17][32]), .s(s[360]), .c_out(c[360]));
    fullAdder fa343 (.a(p[18][30]), .b(p[19][28]), .c_in(p[20][26]), .s(s[361]), .c_out(c[361]));
    fullAdder fa344 (.a(p[21][24]), .b(p[22][22]), .c_in(p[23][20]), .s(s[362]), .c_out(c[362]));
    fullAdder fa345 (.a(p[24][18]), .b(p[25][16]), .c_in(p[26][14]), .s(s[363]), .c_out(c[363]));
    fullAdder fa346 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[07][53]), .c_in(p[08][51]), .s(s[364]), .c_out(c[364]));
    fullAdder fa347 (.a(p[09][49]), .b(p[10][47]), .c_in(p[11][45]), .s(s[365]), .c_out(c[365]));
    fullAdder fa348 (.a(p[12][43]), .b(p[13][41]), .c_in(p[14][39]), .s(s[366]), .c_out(c[366]));
    fullAdder fa349 (.a(p[15][37]), .b(p[16][35]), .c_in(p[17][33]), .s(s[367]), .c_out(c[367]));
    fullAdder fa350 (.a(p[18][31]), .b(p[19][29]), .c_in(mode == 2'b10 ? comp[19] : p[20][27]), .s(s[368]), .c_out(c[368]));
    fullAdder fa351 (.a(p[21][25]), .b(p[22][23]), .c_in(p[23][21]), .s(s[369]), .c_out(c[369]));
    fullAdder fa352 (.a(p[24][19]), .b(p[25][17]), .c_in(p[26][15]), .s(s[370]), .c_out(c[370]));
    fullAdder fa353 (.a(mode == 2'b11 ?  ~comp[07] : 1'b0), .b(p[08][52]), .c_in(p[09][50]), .s(s[371]), .c_out(c[371]));
    fullAdder fa354 (.a(p[10][48]), .b(p[11][46]), .c_in(p[12][44]), .s(s[372]), .c_out(c[372]));
    fullAdder fa355 (.a(p[13][42]), .b(mode == 2'b01 ? comp[14] : p[14][40]), .c_in(p[15][38]), .s(s[373]), .c_out(c[373]));
    fullAdder fa356 (.a(p[16][36]), .b(p[17][34]), .c_in(p[18][32]), .s(s[374]), .c_out(c[374]));
    fullAdder fa357 (.a(p[19][30]), .b(p[20][28]), .c_in(p[21][26]), .s(s[375]), .c_out(c[375]));
    fullAdder fa358 (.a(p[22][24]), .b(p[23][22]), .c_in(p[24][20]), .s(s[376]), .c_out(c[376]));
    halfAdder ha20 (.a(p[25][18]), .b(p[26][16]), .s(s[377]), .c_out(c[377]));
    fullAdder fa359 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[08][53]), .c_in(p[09][51]), .s(s[378]), .c_out(c[378]));
    fullAdder fa360 (.a(p[10][49]), .b(p[11][47]), .c_in(p[12][45]), .s(s[379]), .c_out(c[379]));
    fullAdder fa361 (.a(p[13][43]), .b(mode == 2'b01 ? comp[14] : p[14][41]), .c_in(p[15][39]), .s(s[380]), .c_out(c[380]));
    fullAdder fa362 (.a(p[16][37]), .b(p[17][35]), .c_in(p[18][33]), .s(s[381]), .c_out(c[381]));
    fullAdder fa363 (.a(p[19][31]), .b(p[20][29]), .c_in(mode == 2'b10 ? comp[20] : p[21][27]), .s(s[382]), .c_out(c[382]));
    fullAdder fa364 (.a(p[22][25]), .b(p[23][23]), .c_in(p[24][21]), .s(s[383]), .c_out(c[383]));
    halfAdder ha21 (.a(p[25][19]), .b(p[26][17]), .s(s[384]), .c_out(c[384]));
    fullAdder fa365 (.a(mode == 2'b11 ?  ~comp[08] : 1'b0), .b(p[09][52]), .c_in(p[10][50]), .s(s[385]), .c_out(c[385]));
    fullAdder fa366 (.a(p[11][48]), .b(p[12][46]), .c_in(p[13][44]), .s(s[386]), .c_out(c[386]));
    fullAdder fa367 (.a(mode == 2'b01 ? ~comp[14] : p[14][42]), .b(mode == 2'b01 ? ~comp[15] : p[15][40]), .c_in(p[16][38]), .s(s[387]), .c_out(c[387]));
    fullAdder fa368 (.a(p[17][36]), .b(p[18][34]), .c_in(p[19][32]), .s(s[388]), .c_out(c[388]));
    fullAdder fa369 (.a(p[20][30]), .b(p[21][28]), .c_in(p[22][26]), .s(s[389]), .c_out(c[389]));
    fullAdder fa370 (.a(p[23][24]), .b(p[24][22]), .c_in(p[25][20]), .s(s[390]), .c_out(c[390]));
    fullAdder fa371 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[09][53]), .c_in(p[10][51]), .s(s[391]), .c_out(c[391]));
    fullAdder fa372 (.a(p[11][49]), .b(p[12][47]), .c_in(p[13][45]), .s(s[392]), .c_out(c[392]));
    fullAdder fa373 (.a(p[14][43]), .b(mode == 2'b01 ? 1'b1 : p[15][41]), .c_in(p[16][39]), .s(s[393]), .c_out(c[393]));
    fullAdder fa374 (.a(p[17][37]), .b(p[18][35]), .c_in(p[19][33]), .s(s[394]), .c_out(c[394]));
    fullAdder fa375 (.a(p[20][31]), .b(p[21][29]), .c_in(mode == 2'b10 ? comp[21] : p[22][27]), .s(s[395]), .c_out(c[395]));
    fullAdder fa376 (.a(p[23][25]), .b(p[24][23]), .c_in(p[25][21]), .s(s[396]), .c_out(c[396]));
    fullAdder fa377 (.a(mode == 2'b11 ?  ~comp[09] : 1'b0), .b(p[10][52]), .c_in(p[11][50]), .s(s[397]), .c_out(c[397]));
    fullAdder fa378 (.a(p[12][48]), .b(p[13][46]), .c_in(p[14][44]), .s(s[398]), .c_out(c[398]));
    fullAdder fa379 (.a(p[15][42]), .b(mode == 2'b01 ? ~comp[16] : p[16][40]), .c_in(p[17][38]), .s(s[399]), .c_out(c[399]));
    fullAdder fa380 (.a(p[18][36]), .b(p[19][34]), .c_in(p[20][32]), .s(s[400]), .c_out(c[400]));
    fullAdder fa381 (.a(p[21][30]), .b(p[22][28]), .c_in(p[23][26]), .s(s[401]), .c_out(c[401]));
    fullAdder fa382 (.a(p[24][24]), .b(p[25][22]), .c_in(p[26][20]), .s(s[402]), .c_out(c[402]));
    fullAdder fa383 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[10][53]), .c_in(p[11][51]), .s(s[403]), .c_out(c[403]));
    fullAdder fa384 (.a(p[12][49]), .b(p[13][47]), .c_in(p[14][45]), .s(s[404]), .c_out(c[404]));
    fullAdder fa385 (.a(p[15][43]), .b(mode == 2'b01 ? 1'b1 : p[16][41]), .c_in(p[17][39]), .s(s[405]), .c_out(c[405]));
    fullAdder fa386 (.a(p[18][37]), .b(p[19][35]), .c_in(p[20][33]), .s(s[406]), .c_out(c[406]));
    fullAdder fa387 (.a(p[21][31]), .b(p[22][29]), .c_in(mode == 2'b10 ? comp[22] : p[23][27]), .s(s[407]), .c_out(c[407]));
    fullAdder fa388 (.a(p[24][25]), .b(p[25][23]), .c_in(p[26][21]), .s(s[408]), .c_out(c[408]));
    fullAdder fa389 (.a(mode == 2'b11 ?  ~comp[10] : 1'b0), .b(p[11][52]), .c_in(p[12][50]), .s(s[409]), .c_out(c[409]));
    fullAdder fa390 (.a(p[13][48]), .b(p[14][46]), .c_in(p[15][44]), .s(s[410]), .c_out(c[410]));
    fullAdder fa391 (.a(p[16][42]), .b(mode == 2'b01 ? ~comp[17] : p[17][40]), .c_in(p[18][38]), .s(s[411]), .c_out(c[411]));
    fullAdder fa392 (.a(p[19][36]), .b(p[20][34]), .c_in(p[21][32]), .s(s[412]), .c_out(c[412]));
    fullAdder fa393 (.a(p[22][30]), .b(p[23][28]), .c_in(p[24][26]), .s(s[413]), .c_out(c[413]));
    halfAdder ha22 (.a(p[25][24]), .b(p[26][22]), .s(s[414]), .c_out(c[414]));
    fullAdder fa394 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[11][53]), .c_in(p[12][51]), .s(s[415]), .c_out(c[415]));
    fullAdder fa395 (.a(p[13][49]), .b(p[14][47]), .c_in(p[15][45]), .s(s[416]), .c_out(c[416]));
    fullAdder fa396 (.a(p[16][43]), .b(mode == 2'b01 ? 1'b1 : p[17][41]), .c_in(p[18][39]), .s(s[417]), .c_out(c[417]));
    fullAdder fa397 (.a(p[19][37]), .b(p[20][35]), .c_in(p[21][33]), .s(s[418]), .c_out(c[418]));
    fullAdder fa398 (.a(p[22][31]), .b(p[23][29]), .c_in(mode == 2'b10 ? comp[23] : p[24][27]), .s(s[419]), .c_out(c[419]));
    halfAdder ha23 (.a(p[25][25]), .b(p[26][23]), .s(s[420]), .c_out(c[420]));
    fullAdder fa399 (.a(mode == 2'b11 ?  ~comp[11] : 1'b0), .b(p[12][52]), .c_in(p[13][50]), .s(s[421]), .c_out(c[421]));
    fullAdder fa400 (.a(p[14][48]), .b(p[15][46]), .c_in(p[16][44]), .s(s[422]), .c_out(c[422]));
    fullAdder fa401 (.a(p[17][42]), .b(mode == 2'b01 ? ~comp[18] : p[18][40]), .c_in(p[19][38]), .s(s[423]), .c_out(c[423]));
    fullAdder fa402 (.a(p[20][36]), .b(p[21][34]), .c_in(p[22][32]), .s(s[424]), .c_out(c[424]));
    fullAdder fa403 (.a(p[23][30]), .b(p[24][28]), .c_in(p[25][26]), .s(s[425]), .c_out(c[425]));
    fullAdder fa404 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[12][53]), .c_in(p[13][51]), .s(s[426]), .c_out(c[426]));
    fullAdder fa405 (.a(p[14][49]), .b(p[15][47]), .c_in(p[16][45]), .s(s[427]), .c_out(c[427]));
    fullAdder fa406 (.a(p[17][43]), .b(mode == 2'b01 ? 1'b1 : p[18][41]), .c_in(p[19][39]), .s(s[428]), .c_out(c[428]));
    fullAdder fa407 (.a(p[20][37]), .b(p[21][35]), .c_in(p[22][33]), .s(s[429]), .c_out(c[429]));
    fullAdder fa408 (.a(p[23][31]), .b(p[24][29]), .c_in(mode == 2'b10 ? comp[24] : p[25][27]), .s(s[430]), .c_out(c[430]));
    fullAdder fa409 (.a(mode == 2'b11 ?  ~comp[12] : 1'b0), .b(p[13][52]), .c_in(p[14][50]), .s(s[431]), .c_out(c[431]));
    fullAdder fa410 (.a(p[15][48]), .b(p[16][46]), .c_in(p[17][44]), .s(s[432]), .c_out(c[432]));
    fullAdder fa411 (.a(p[18][42]), .b(p[19][40]), .c_in(p[20][38]), .s(s[433]), .c_out(c[433]));
    fullAdder fa412 (.a(p[21][36]), .b(p[22][34]), .c_in(p[23][32]), .s(s[434]), .c_out(c[434]));
    fullAdder fa413 (.a(p[24][30]), .b(p[25][28]), .c_in(p[26][26]), .s(s[435]), .c_out(c[435]));
    fullAdder fa414 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[13][53]), .c_in(p[14][51]), .s(s[436]), .c_out(c[436]));
    fullAdder fa415 (.a(p[15][49]), .b(p[16][47]), .c_in(p[17][45]), .s(s[437]), .c_out(c[437]));
    fullAdder fa416 (.a(p[18][43]), .b(p[19][41]), .c_in(p[20][39]), .s(s[438]), .c_out(c[438]));
    fullAdder fa417 (.a(p[21][37]), .b(p[22][35]), .c_in(p[23][33]), .s(s[439]), .c_out(c[439]));
    fullAdder fa418 (.a(p[24][31]), .b(p[25][29]), .c_in(mode == 2'b10 ? comp[25] : p[26][27]), .s(s[440]), .c_out(c[440]));
    fullAdder fa419 (.a(mode == 2'b11 ?  ~comp[13] : 1'b0), .b(p[14][52]), .c_in(p[15][50]), .s(s[441]), .c_out(c[441]));
    fullAdder fa420 (.a(p[16][48]), .b(p[17][46]), .c_in(p[18][44]), .s(s[442]), .c_out(c[442]));
    fullAdder fa421 (.a(p[19][42]), .b(p[20][40]), .c_in(p[21][38]), .s(s[443]), .c_out(c[443]));
    fullAdder fa422 (.a(p[22][36]), .b(p[23][34]), .c_in(p[24][32]), .s(s[444]), .c_out(c[444]));
    halfAdder ha24 (.a(p[25][30]), .b(p[26][28]), .s(s[445]), .c_out(c[445]));
    fullAdder fa423 (.a(mode == 2'b11 ? 1'b1 : 1'b0), .b(p[14][53]), .c_in(p[15][51]), .s(s[446]), .c_out(c[446]));
    fullAdder fa424 (.a(p[16][49]), .b(p[17][47]), .c_in(p[18][45]), .s(s[447]), .c_out(c[447]));
    fullAdder fa425 (.a(p[19][43]), .b(p[20][41]), .c_in(p[21][39]), .s(s[448]), .c_out(c[448]));
    fullAdder fa426 (.a(p[22][37]), .b(p[23][35]), .c_in(p[24][33]), .s(s[449]), .c_out(c[449]));
    halfAdder ha25 (.a(p[25][31]), .b(p[26][29]), .s(s[450]), .c_out(c[450]));
    fullAdder fa427 (.a(mode == 2'b11 ?  ~comp[14] : mode == 2'b10 ?  comp[14] : 1'b0), .b(p[15][52]), .c_in(p[16][50]), .s(s[451]), .c_out(c[451]));
    fullAdder fa428 (.a(p[17][48]), .b(p[18][46]), .c_in(p[19][44]), .s(s[452]), .c_out(c[452]));
    fullAdder fa429 (.a(p[20][42]), .b(p[21][40]), .c_in(p[22][38]), .s(s[453]), .c_out(c[453]));
    fullAdder fa430 (.a(p[23][36]), .b(p[24][34]), .c_in(p[25][32]), .s(s[454]), .c_out(c[454]));
    fullAdder fa431 (.a(mode == 2'b11 ?  1'b1 : mode == 2'b10 ?  comp[14] : 1'b0), .b(p[15][53]), .c_in(p[16][51]), .s(s[455]), .c_out(c[455]));
    fullAdder fa432 (.a(p[17][49]), .b(p[18][47]), .c_in(p[19][45]), .s(s[456]), .c_out(c[456]));
    fullAdder fa433 (.a(p[20][43]), .b(p[21][41]), .c_in(p[22][39]), .s(s[457]), .c_out(c[457]));
    fullAdder fa434 (.a(p[23][37]), .b(p[24][35]), .c_in(p[25][33]), .s(s[458]), .c_out(c[458]));
    fullAdder fa435 (.a(mode == 2'b10 ?  ~comp[14] : 1'b0), .b(mode[1] == 1'b1 ?  ~comp[15] : 1'b0), .c_in(p[16][52]), .s(s[459]), .c_out(c[459]));
    fullAdder fa436 (.a(p[17][50]), .b(p[18][48]), .c_in(p[19][46]), .s(s[460]), .c_out(c[460]));
    fullAdder fa437 (.a(p[20][44]), .b(p[21][42]), .c_in(mode == 2'b01 ? comp[21] : p[22][40]), .s(s[461]), .c_out(c[461]));
    fullAdder fa438 (.a(p[23][38]), .b(p[24][36]), .c_in(p[25][34]), .s(s[462]), .c_out(c[462]));
    fullAdder fa439 (.a(mode[1] == 1'b1 ? 1'b1 : 1'b0), .b(p[16][53]), .c_in(p[17][51]), .s(s[463]), .c_out(c[463]));
    fullAdder fa440 (.a(p[18][49]), .b(p[19][47]), .c_in(p[20][45]), .s(s[464]), .c_out(c[464]));
    fullAdder fa441 (.a(p[21][43]), .b(p[22][41]), .c_in(p[23][39]), .s(s[465]), .c_out(c[465]));
    fullAdder fa442 (.a(p[24][37]), .b(p[25][35]), .c_in(p[26][33]), .s(s[466]), .c_out(c[466]));
    fullAdder fa443 (.a(mode[1] == 1'b1 ? ~comp[16] : 1'b0), .b(p[17][52]), .c_in(p[18][50]), .s(s[467]), .c_out(c[467]));
    fullAdder fa444 (.a(p[19][48]), .b(p[20][46]), .c_in(p[21][44]), .s(s[468]), .c_out(c[468]));
    fullAdder fa445 (.a(p[22][42]), .b(mode == 2'b01 ? comp[22] : p[23][40]), .c_in(p[24][38]), .s(s[469]), .c_out(c[469]));
    halfAdder ha26 (.a(p[25][36]), .b(p[26][34]), .s(s[470]), .c_out(c[470]));
    fullAdder fa446 (.a(mode[1] == 1'b1 ? 1'b1: 1'b0), .b(p[17][53]), .c_in(p[18][51]), .s(s[471]), .c_out(c[471]));
    fullAdder fa447 (.a(p[19][49]), .b(p[20][47]), .c_in(p[21][45]), .s(s[472]), .c_out(c[472]));
    fullAdder fa448 (.a(p[22][43]), .b(p[23][41]), .c_in(p[24][39]), .s(s[473]), .c_out(c[473]));
    halfAdder ha27 (.a(p[25][37]), .b(p[26][35]), .s(s[474]), .c_out(c[474]));
    fullAdder fa449 (.a(mode[1] == 1'b1 ? ~comp[17] : 1'b0), .b(p[18][52]), .c_in(p[19][50]), .s(s[475]), .c_out(c[475]));
    fullAdder fa450 (.a(p[20][48]), .b(p[21][46]), .c_in(p[22][44]), .s(s[476]), .c_out(c[476]));
    fullAdder fa451 (.a(p[23][42]), .b(mode == 2'b01 ? comp[23] : p[24][40]), .c_in(p[25][38]), .s(s[477]), .c_out(c[477]));
    fullAdder fa452 (.a(mode[1] == 1'b1 ? 1'b1 : 1'b0), .b(p[18][53]), .c_in(p[19][51]), .s(s[478]), .c_out(c[478]));
    fullAdder fa453 (.a(p[20][49]), .b(p[21][47]), .c_in(p[22][45]), .s(s[479]), .c_out(c[479]));
    fullAdder fa454 (.a(p[23][43]), .b(p[24][41]), .c_in(p[25][39]), .s(s[480]), .c_out(c[480]));
    fullAdder fa455 (.a(mode[1] == 1'b1 ? ~comp[18] : 1'b0), .b(p[19][52]), .c_in(p[20][50]), .s(s[481]), .c_out(c[481]));
    fullAdder fa456 (.a(p[21][48]), .b(p[22][46]), .c_in(p[23][44]), .s(s[482]), .c_out(c[482]));
    fullAdder fa457 (.a(p[24][42]), .b(mode == 2'b01 ? comp[24] : p[25][40]), .c_in(p[26][38]), .s(s[483]), .c_out(c[483]));
    fullAdder fa458 (.a(mode[1] == 1'b1 ? 1'b1 : 1'b0), .b(p[19][53]), .c_in(p[20][51]), .s(s[484]), .c_out(c[484]));
    fullAdder fa459 (.a(p[21][49]), .b(p[22][47]), .c_in(p[23][45]), .s(s[485]), .c_out(c[485]));
    fullAdder fa460 (.a(p[24][43]), .b(p[25][41]), .c_in(p[26][39]), .s(s[486]), .c_out(c[486]));
    fullAdder fa461 (.a(mode[1] == 1'b1 ? ~comp[19] : 1'b0), .b(p[20][52]), .c_in(p[21][50]), .s(s[487]), .c_out(c[487]));
    fullAdder fa462 (.a(p[22][48]), .b(p[23][46]), .c_in(p[24][44]), .s(s[488]), .c_out(c[488]));
    halfAdder ha28 (.a(p[25][42]), .b(mode == 2'b01 ? comp[25] : p[26][40]), .s(s[489]), .c_out(c[489]));
    fullAdder fa463 (.a(mode[1] == 1'b1 ? 1'b1 : 1'b0), .b(p[20][53]), .c_in(p[21][51]), .s(s[490]), .c_out(c[490]));
    fullAdder fa464 (.a(p[22][49]), .b(p[23][47]), .c_in(p[24][45]), .s(s[491]), .c_out(c[491]));
    halfAdder ha29 (.a(p[25][43]), .b(p[26][41]), .s(s[492]), .c_out(c[492]));
    fullAdder fa465 (.a(mode[1] == 1'b1 ? ~comp[20] : 1'b0), .b(p[21][52]), .c_in(p[22][50]), .s(s[493]), .c_out(c[493]));
    fullAdder fa466 (.a(p[23][48]), .b(p[24][46]), .c_in(p[25][44]), .s(s[494]), .c_out(c[494]));
    fullAdder fa467 (.a(mode[1] == 1'b1 ? 1'b1 : 1'b0), .b(p[21][53]), .c_in(p[22][51]), .s(s[495]), .c_out(c[495]));
    fullAdder fa468 (.a(p[23][49]), .b(p[24][47]), .c_in(p[25][45]), .s(s[496]), .c_out(c[496]));
    fullAdder fa469 (.a(mode[1] == 1'b1 ? ~comp[21] : mode[0] ==1'b1 ? comp[21] : 1'b0), .b(p[22][52]), .c_in(p[23][50]), .s(s[497]), .c_out(c[497]));
    fullAdder fa470 (.a(p[24][48]), .b(p[25][46]), .c_in(p[26][44]), .s(s[498]), .c_out(c[498]));
    fullAdder fa471 (.a(mode[1] == 1'b1 ? 1'b1 :  mode[0] ==1'b1 ? comp[21] : 1'b0), .b(p[22][53]), .c_in(p[23][51]), .s(s[499]), .c_out(c[499]));
    fullAdder fa472 (.a(p[24][49]), .b(p[25][47]), .c_in(p[26][45]), .s(s[500]), .c_out(c[500]));
    fullAdder fa473 (.a(mode ==  2'b01 ? ~comp[21] :1'b0), .b(~comp[22]), .c_in(p[23][52]), .s(s[501]), .c_out(c[501]));
    fullAdder fa474 (.a(p[24][50]), .b(p[25][48]), .c_in(p[26][46]), .s(s[502]), .c_out(c[502]));
    fullAdder fa475 (.a(1'b1), .b(p[23][53]), .c_in(p[24][51]), .s(s[503]), .c_out(c[503]));
    halfAdder ha30 (.a(p[25][49]), .b(p[26][47]), .s(s[504]), .c_out(c[504]));
    fullAdder fa476 (.a(~comp[23]), .b(p[24][52]), .c_in(p[25][50]), .s(s[505]), .c_out(c[505]));
    fullAdder fa477 (.a(1'b1), .b(p[24][53]), .c_in(p[25][51]), .s(s[506]), .c_out(c[506]));
    fullAdder fa478 (.a(~comp[24]), .b(p[25][52]), .c_in(p[26][50]), .s(s[507]), .c_out(c[507]));
    fullAdder fa479 (.a(1'b1), .b(p[25][53]), .c_in(p[26][51]), .s(s[508]), .c_out(c[508]));
    // Stage 2 Reduction
    fullAdder fa480 (.a(p[00][03]), .b(c[0]), .c_in(p[01][01]), .s(s[509]), .c_out(c[509]));
    fullAdder fa481 (.a(s[3]), .b(c[2]), .c_in(s[4]), .s(s[510]), .c_out(c[510]));
    fullAdder fa482 (.a(s[5]), .b(c[3]), .c_in(p[03][01]), .s(s[511]), .c_out(c[511]));
    fullAdder fa483 (.a(s[6]), .b(c[5]), .c_in(s[7]), .s(s[512]), .c_out(c[512]));
    fullAdder fa484 (.a(s[8]), .b(c[6]), .c_in(s[9]), .s(s[513]), .c_out(c[513]));
    fullAdder fa485 (.a(s[10]), .b(c[8]), .c_in(s[11]), .s(s[514]), .c_out(c[514]));
    halfAdder ha31 (.a(c[9]), .b(mode == 2'b01 ? 1'b0 : comp[5]), .s(s[515]), .c_out(c[515]));
    fullAdder fa486 (.a(s[12]), .b(c[10]), .c_in(s[13]), .s(s[516]), .c_out(c[516]));
    fullAdder fa487 (.a(s[14]), .b(c[12]), .c_in(s[15]), .s(s[517]), .c_out(c[517]));
    halfAdder ha32 (.a(c[13]), .b(s[16]), .s(s[518]), .c_out(c[518]));
    fullAdder fa488 (.a(s[17]), .b(c[14]), .c_in(s[18]), .s(s[519]), .c_out(c[519]));
    fullAdder fa489 (.a(c[15]), .b(p[06][01]), .c_in(c[16]), .s(s[520]), .c_out(c[520]));
    fullAdder fa490 (.a(s[19]), .b(c[17]), .c_in(s[20]), .s(s[521]), .c_out(c[521]));
    halfAdder ha33 (.a(c[18]), .b(s[21]), .s(s[522]), .c_out(c[522]));
    fullAdder fa491 (.a(s[22]), .b(c[19]), .c_in(s[23]), .s(s[523]), .c_out(c[523]));
    fullAdder fa492 (.a(c[20]), .b(s[24]), .c_in(c[21]), .s(s[524]), .c_out(c[524]));
    fullAdder fa493 (.a(s[25]), .b(c[22]), .c_in(s[26]), .s(s[525]), .c_out(c[525]));
    fullAdder fa494 (.a(c[23]), .b(s[27]), .c_in(c[24]), .s(s[526]), .c_out(c[526]));
    fullAdder fa495 (.a(s[28]), .b(c[25]), .c_in(s[29]), .s(s[527]), .c_out(c[527]));
    fullAdder fa496 (.a(c[26]), .b(s[30]), .c_in(c[27]), .s(s[528]), .c_out(c[528]));
    fullAdder fa497 (.a(s[31]), .b(c[28]), .c_in(s[32]), .s(s[529]), .c_out(c[529]));
    fullAdder fa498 (.a(c[29]), .b(s[33]), .c_in(c[30]), .s(s[530]), .c_out(c[530]));
    fullAdder fa499 (.a(s[35]), .b(c[31]), .c_in(s[36]), .s(s[531]), .c_out(c[531]));
    fullAdder fa500 (.a(c[32]), .b(s[37]), .c_in(c[33]), .s(s[532]), .c_out(c[532]));
    halfAdder ha34 (.a(p[09][01]), .b(c[34]), .s(s[533]), .c_out(c[533]));
    fullAdder fa501 (.a(s[38]), .b(c[35]), .c_in(s[39]), .s(s[534]), .c_out(c[534]));
    fullAdder fa502 (.a(c[36]), .b(s[40]), .c_in(c[37]), .s(s[535]), .c_out(c[535]));
    fullAdder fa503 (.a(s[42]), .b(c[38]), .c_in(s[43]), .s(s[536]), .c_out(c[536]));
    fullAdder fa504 (.a(c[39]), .b(s[44]), .c_in(c[40]), .s(s[537]), .c_out(c[537]));
    halfAdder ha35 (.a(s[45]), .b(c[41]), .s(s[538]), .c_out(c[538]));
    fullAdder fa505 (.a(s[46]), .b(c[42]), .c_in(s[47]), .s(s[539]), .c_out(c[539]));
    fullAdder fa506 (.a(c[43]), .b(s[48]), .c_in(c[44]), .s(s[540]), .c_out(c[540]));
    fullAdder fa507 (.a(s[49]), .b(c[45]), .c_in(mode == 2'b01 ? 1'b0 : comp[11]), .s(s[541]), .c_out(c[541]));
    fullAdder fa508 (.a(s[50]), .b(c[46]), .c_in(s[51]), .s(s[542]), .c_out(c[542]));
    fullAdder fa509 (.a(c[47]), .b(s[52]), .c_in(c[48]), .s(s[543]), .c_out(c[543]));
    halfAdder ha36 (.a(s[53]), .b(c[49]), .s(s[544]), .c_out(c[544]));
    fullAdder fa510 (.a(s[54]), .b(c[50]), .c_in(s[55]), .s(s[545]), .c_out(c[545]));
    fullAdder fa511 (.a(c[51]), .b(s[56]), .c_in(c[52]), .s(s[546]), .c_out(c[546]));
    fullAdder fa512 (.a(s[57]), .b(c[53]), .c_in(s[58]), .s(s[547]), .c_out(c[547]));
    fullAdder fa513 (.a(s[59]), .b(c[54]), .c_in(s[60]), .s(s[548]), .c_out(c[548]));
    fullAdder fa514 (.a(c[55]), .b(s[61]), .c_in(c[56]), .s(s[549]), .c_out(c[549]));
    fullAdder fa515 (.a(s[62]), .b(c[57]), .c_in(p[12][01]), .s(s[550]), .c_out(c[550]));
    fullAdder fa516 (.a(s[63]), .b(c[59]), .c_in(s[64]), .s(s[551]), .c_out(c[551]));
    fullAdder fa517 (.a(c[60]), .b(s[65]), .c_in(c[61]), .s(s[552]), .c_out(c[552]));
    fullAdder fa518 (.a(s[66]), .b(c[62]), .c_in(s[67]), .s(s[553]), .c_out(c[553]));
    fullAdder fa519 (.a(s[68]), .b(c[63]), .c_in(s[69]), .s(s[554]), .c_out(c[554]));
    fullAdder fa520 (.a(c[64]), .b(s[70]), .c_in(c[65]), .s(s[555]), .c_out(c[555]));
    fullAdder fa521 (.a(s[71]), .b(c[66]), .c_in(s[72]), .s(s[556]), .c_out(c[556]));
    fullAdder fa522 (.a(s[73]), .b(c[68]), .c_in(s[74]), .s(s[557]), .c_out(c[557]));
    fullAdder fa523 (.a(c[69]), .b(s[75]), .c_in(c[70]), .s(s[558]), .c_out(c[558]));
    fullAdder fa524 (.a(s[76]), .b(c[71]), .c_in(s[77]), .s(s[559]), .c_out(c[559]));
    halfAdder ha37 (.a(c[72]), .b(mode == 2'b11 ? comp[14] : 1'b0), .s(s[560]), .c_out(c[560]));
    fullAdder fa525 (.a(s[78]), .b(c[73]), .c_in(s[79]), .s(s[561]), .c_out(c[561]));
    fullAdder fa526 (.a(c[74]), .b(s[80]), .c_in(c[75]), .s(s[562]), .c_out(c[562]));
    fullAdder fa527 (.a(s[81]), .b(c[76]), .c_in(s[82]), .s(s[563]), .c_out(c[563]));
    fullAdder fa528 (.a(s[83]), .b(c[78]), .c_in(s[84]), .s(s[564]), .c_out(c[564]));
    fullAdder fa529 (.a(c[79]), .b(s[85]), .c_in(c[80]), .s(s[565]), .c_out(c[565]));
    fullAdder fa530 (.a(s[86]), .b(c[81]), .c_in(s[87]), .s(s[566]), .c_out(c[566]));
    halfAdder ha38 (.a(c[82]), .b(s[88]), .s(s[567]), .c_out(c[567]));
    fullAdder fa531 (.a(s[89]), .b(c[83]), .c_in(s[90]), .s(s[568]), .c_out(c[568]));
    fullAdder fa532 (.a(c[84]), .b(s[91]), .c_in(c[85]), .s(s[569]), .c_out(c[569]));
    fullAdder fa533 (.a(s[92]), .b(c[86]), .c_in(s[93]), .s(s[570]), .c_out(c[570]));
    fullAdder fa534 (.a(c[87]), .b(p[15][01]), .c_in(c[88]), .s(s[571]), .c_out(c[571]));
    fullAdder fa535 (.a(s[94]), .b(c[89]), .c_in(s[95]), .s(s[572]), .c_out(c[572]));
    fullAdder fa536 (.a(c[90]), .b(s[96]), .c_in(c[91]), .s(s[573]), .c_out(c[573]));
    fullAdder fa537 (.a(s[97]), .b(c[92]), .c_in(s[98]), .s(s[574]), .c_out(c[574]));
    halfAdder ha39 (.a(c[93]), .b(s[99]), .s(s[575]), .c_out(c[575]));
    fullAdder fa538 (.a(s[100]), .b(c[94]), .c_in(s[101]), .s(s[576]), .c_out(c[576]));
    fullAdder fa539 (.a(c[95]), .b(s[102]), .c_in(c[96]), .s(s[577]), .c_out(c[577]));
    fullAdder fa540 (.a(s[103]), .b(c[97]), .c_in(s[104]), .s(s[578]), .c_out(c[578]));
    fullAdder fa541 (.a(c[98]), .b(s[105]), .c_in(c[99]), .s(s[579]), .c_out(c[579]));
    fullAdder fa542 (.a(s[106]), .b(c[100]), .c_in(s[107]), .s(s[580]), .c_out(c[580]));
    fullAdder fa543 (.a(c[101]), .b(s[108]), .c_in(c[102]), .s(s[581]), .c_out(c[581]));
    fullAdder fa544 (.a(s[109]), .b(c[103]), .c_in(s[110]), .s(s[582]), .c_out(c[582]));
    fullAdder fa545 (.a(c[104]), .b(s[111]), .c_in(c[105]), .s(s[583]), .c_out(c[583]));
    fullAdder fa546 (.a(s[112]), .b(c[106]), .c_in(s[113]), .s(s[584]), .c_out(c[584]));
    fullAdder fa547 (.a(c[107]), .b(s[114]), .c_in(c[108]), .s(s[585]), .c_out(c[585]));
    fullAdder fa548 (.a(s[115]), .b(c[109]), .c_in(s[116]), .s(s[586]), .c_out(c[586]));
    fullAdder fa549 (.a(c[110]), .b(s[117]), .c_in(c[111]), .s(s[587]), .c_out(c[587]));
    fullAdder fa550 (.a(s[118]), .b(c[112]), .c_in(s[119]), .s(s[588]), .c_out(c[588]));
    fullAdder fa551 (.a(c[113]), .b(s[120]), .c_in(c[114]), .s(s[589]), .c_out(c[589]));
    fullAdder fa552 (.a(s[121]), .b(c[115]), .c_in(s[122]), .s(s[590]), .c_out(c[590]));
    fullAdder fa553 (.a(c[116]), .b(s[123]), .c_in(c[117]), .s(s[591]), .c_out(c[591]));
    fullAdder fa554 (.a(s[125]), .b(c[118]), .c_in(s[126]), .s(s[592]), .c_out(c[592]));
    fullAdder fa555 (.a(c[119]), .b(s[127]), .c_in(c[120]), .s(s[593]), .c_out(c[593]));
    fullAdder fa556 (.a(s[128]), .b(c[121]), .c_in(s[129]), .s(s[594]), .c_out(c[594]));
    fullAdder fa557 (.a(c[122]), .b(s[130]), .c_in(c[123]), .s(s[595]), .c_out(c[595]));
    halfAdder ha40 (.a(p[18][01]), .b(c[124]), .s(s[596]), .c_out(c[596]));
    fullAdder fa558 (.a(s[131]), .b(c[125]), .c_in(s[132]), .s(s[597]), .c_out(c[597]));
    fullAdder fa559 (.a(c[126]), .b(s[133]), .c_in(c[127]), .s(s[598]), .c_out(c[598]));
    fullAdder fa560 (.a(s[134]), .b(c[128]), .c_in(s[135]), .s(s[599]), .c_out(c[599]));
    fullAdder fa561 (.a(c[129]), .b(s[136]), .c_in(c[130]), .s(s[600]), .c_out(c[600]));
    fullAdder fa562 (.a(s[138]), .b(c[131]), .c_in(s[139]), .s(s[601]), .c_out(c[601]));
    fullAdder fa563 (.a(c[132]), .b(s[140]), .c_in(c[133]), .s(s[602]), .c_out(c[602]));
    fullAdder fa564 (.a(s[141]), .b(c[134]), .c_in(s[142]), .s(s[603]), .c_out(c[603]));
    fullAdder fa565 (.a(c[135]), .b(s[143]), .c_in(c[136]), .s(s[604]), .c_out(c[604]));
    halfAdder ha41 (.a(s[144]), .b(c[137]), .s(s[605]), .c_out(c[605]));
    fullAdder fa566 (.a(s[145]), .b(c[138]), .c_in(s[146]), .s(s[606]), .c_out(c[606]));
    fullAdder fa567 (.a(c[139]), .b(s[147]), .c_in(c[140]), .s(s[607]), .c_out(c[607]));
    fullAdder fa568 (.a(s[148]), .b(c[141]), .c_in(s[149]), .s(s[608]), .c_out(c[608]));
    fullAdder fa569 (.a(c[142]), .b(s[150]), .c_in(c[143]), .s(s[609]), .c_out(c[609]));
    fullAdder fa570 (.a(s[151]), .b(c[144]), .c_in(mode == 2'b11 ? comp[20] : 1'b0), .s(s[610]), .c_out(c[610]));
    fullAdder fa571 (.a(s[152]), .b(c[145]), .c_in(s[153]), .s(s[611]), .c_out(c[611]));
    fullAdder fa572 (.a(c[146]), .b(s[154]), .c_in(c[147]), .s(s[612]), .c_out(c[612]));
    fullAdder fa573 (.a(s[155]), .b(c[148]), .c_in(s[156]), .s(s[613]), .c_out(c[613]));
    fullAdder fa574 (.a(c[149]), .b(s[157]), .c_in(c[150]), .s(s[614]), .c_out(c[614]));
    halfAdder ha42 (.a(s[158]), .b(c[151]), .s(s[615]), .c_out(c[615]));
    fullAdder fa575 (.a(s[159]), .b(c[152]), .c_in(s[160]), .s(s[616]), .c_out(c[616]));
    fullAdder fa576 (.a(c[153]), .b(s[161]), .c_in(c[154]), .s(s[617]), .c_out(c[617]));
    fullAdder fa577 (.a(s[162]), .b(c[155]), .c_in(s[163]), .s(s[618]), .c_out(c[618]));
    fullAdder fa578 (.a(c[156]), .b(s[164]), .c_in(c[157]), .s(s[619]), .c_out(c[619]));
    fullAdder fa579 (.a(s[165]), .b(c[158]), .c_in(s[166]), .s(s[620]), .c_out(c[620]));
    fullAdder fa580 (.a(s[167]), .b(c[159]), .c_in(s[168]), .s(s[621]), .c_out(c[621]));
    fullAdder fa581 (.a(c[160]), .b(s[169]), .c_in(c[161]), .s(s[622]), .c_out(c[622]));
    fullAdder fa582 (.a(s[170]), .b(c[162]), .c_in(s[171]), .s(s[623]), .c_out(c[623]));
    fullAdder fa583 (.a(c[163]), .b(s[172]), .c_in(c[164]), .s(s[624]), .c_out(c[624]));
    fullAdder fa584 (.a(s[173]), .b(c[165]), .c_in(p[21][01]), .s(s[625]), .c_out(c[625]));
    fullAdder fa585 (.a(s[174]), .b(c[167]), .c_in(s[175]), .s(s[626]), .c_out(c[626]));
    fullAdder fa586 (.a(c[168]), .b(s[176]), .c_in(c[169]), .s(s[627]), .c_out(c[627]));
    fullAdder fa587 (.a(s[177]), .b(c[170]), .c_in(s[178]), .s(s[628]), .c_out(c[628]));
    fullAdder fa588 (.a(c[171]), .b(s[179]), .c_in(c[172]), .s(s[629]), .c_out(c[629]));
    fullAdder fa589 (.a(s[180]), .b(c[173]), .c_in(s[181]), .s(s[630]), .c_out(c[630]));
    fullAdder fa590 (.a(s[182]), .b(c[174]), .c_in(s[183]), .s(s[631]), .c_out(c[631]));
    fullAdder fa591 (.a(c[175]), .b(s[184]), .c_in(c[176]), .s(s[632]), .c_out(c[632]));
    fullAdder fa592 (.a(s[185]), .b(c[177]), .c_in(s[186]), .s(s[633]), .c_out(c[633]));
    fullAdder fa593 (.a(c[178]), .b(s[187]), .c_in(c[179]), .s(s[634]), .c_out(c[634]));
    fullAdder fa594 (.a(s[188]), .b(c[180]), .c_in(s[189]), .s(s[635]), .c_out(c[635]));
    fullAdder fa595 (.a(s[190]), .b(c[182]), .c_in(s[191]), .s(s[636]), .c_out(c[636]));
    fullAdder fa596 (.a(c[183]), .b(s[192]), .c_in(c[184]), .s(s[637]), .c_out(c[637]));
    fullAdder fa597 (.a(s[193]), .b(c[185]), .c_in(s[194]), .s(s[638]), .c_out(c[638]));
    fullAdder fa598 (.a(c[186]), .b(s[195]), .c_in(c[187]), .s(s[639]), .c_out(c[639]));
    fullAdder fa599 (.a(s[196]), .b(c[188]), .c_in(s[197]), .s(s[640]), .c_out(c[640]));
    halfAdder ha43 (.a(c[189]), .b(mode == 2'b11 ? comp[23] : 1'b0), .s(s[641]), .c_out(c[641]));
    fullAdder fa600 (.a(s[198]), .b(c[190]), .c_in(s[199]), .s(s[642]), .c_out(c[642]));
    fullAdder fa601 (.a(c[191]), .b(s[200]), .c_in(c[192]), .s(s[643]), .c_out(c[643]));
    fullAdder fa602 (.a(s[201]), .b(c[193]), .c_in(s[202]), .s(s[644]), .c_out(c[644]));
    fullAdder fa603 (.a(c[194]), .b(s[203]), .c_in(c[195]), .s(s[645]), .c_out(c[645]));
    fullAdder fa604 (.a(s[204]), .b(c[196]), .c_in(s[205]), .s(s[646]), .c_out(c[646]));
    fullAdder fa605 (.a(s[206]), .b(c[198]), .c_in(s[207]), .s(s[647]), .c_out(c[647]));
    fullAdder fa606 (.a(c[199]), .b(s[208]), .c_in(c[200]), .s(s[648]), .c_out(c[648]));
    fullAdder fa607 (.a(s[209]), .b(c[201]), .c_in(s[210]), .s(s[649]), .c_out(c[649]));
    fullAdder fa608 (.a(c[202]), .b(s[211]), .c_in(c[203]), .s(s[650]), .c_out(c[650]));
    fullAdder fa609 (.a(s[212]), .b(c[204]), .c_in(s[213]), .s(s[651]), .c_out(c[651]));
    halfAdder ha44 (.a(c[205]), .b(s[214]), .s(s[652]), .c_out(c[652]));
    fullAdder fa610 (.a(s[215]), .b(c[206]), .c_in(s[216]), .s(s[653]), .c_out(c[653]));
    fullAdder fa611 (.a(c[207]), .b(s[217]), .c_in(c[208]), .s(s[654]), .c_out(c[654]));
    fullAdder fa612 (.a(s[218]), .b(c[209]), .c_in(s[219]), .s(s[655]), .c_out(c[655]));
    fullAdder fa613 (.a(c[210]), .b(s[220]), .c_in(c[211]), .s(s[656]), .c_out(c[656]));
    fullAdder fa614 (.a(s[221]), .b(c[212]), .c_in(s[222]), .s(s[657]), .c_out(c[657]));
    fullAdder fa615 (.a(c[213]), .b(p[24][01]), .c_in(c[214]), .s(s[658]), .c_out(c[658]));
    fullAdder fa616 (.a(s[223]), .b(c[215]), .c_in(s[224]), .s(s[659]), .c_out(c[659]));
    fullAdder fa617 (.a(c[216]), .b(s[225]), .c_in(c[217]), .s(s[660]), .c_out(c[660]));
    fullAdder fa618 (.a(s[226]), .b(c[218]), .c_in(s[227]), .s(s[661]), .c_out(c[661]));
    fullAdder fa619 (.a(c[219]), .b(s[228]), .c_in(c[220]), .s(s[662]), .c_out(c[662]));
    fullAdder fa620 (.a(s[229]), .b(c[221]), .c_in(s[230]), .s(s[663]), .c_out(c[663]));
    halfAdder ha45 (.a(c[222]), .b(s[231]), .s(s[664]), .c_out(c[664]));
    fullAdder fa621 (.a(s[232]), .b(c[223]), .c_in(s[233]), .s(s[665]), .c_out(c[665]));
    fullAdder fa622 (.a(c[224]), .b(s[234]), .c_in(c[225]), .s(s[666]), .c_out(c[666]));
    fullAdder fa623 (.a(s[235]), .b(c[226]), .c_in(s[236]), .s(s[667]), .c_out(c[667]));
    fullAdder fa624 (.a(c[227]), .b(s[237]), .c_in(c[228]), .s(s[668]), .c_out(c[668]));
    fullAdder fa625 (.a(s[238]), .b(c[229]), .c_in(s[239]), .s(s[669]), .c_out(c[669]));
    fullAdder fa626 (.a(c[230]), .b(s[240]), .c_in(c[231]), .s(s[670]), .c_out(c[670]));
    fullAdder fa627 (.a(s[241]), .b(c[232]), .c_in(s[242]), .s(s[671]), .c_out(c[671]));
    fullAdder fa628 (.a(c[233]), .b(s[243]), .c_in(c[234]), .s(s[672]), .c_out(c[672]));
    fullAdder fa629 (.a(s[244]), .b(c[235]), .c_in(s[245]), .s(s[673]), .c_out(c[673]));
    fullAdder fa630 (.a(c[236]), .b(s[246]), .c_in(c[237]), .s(s[674]), .c_out(c[674]));
    fullAdder fa631 (.a(s[247]), .b(c[238]), .c_in(s[248]), .s(s[675]), .c_out(c[675]));
    fullAdder fa632 (.a(c[239]), .b(s[249]), .c_in(c[240]), .s(s[676]), .c_out(c[676]));
    fullAdder fa633 (.a(s[250]), .b(c[241]), .c_in(s[251]), .s(s[677]), .c_out(c[677]));
    fullAdder fa634 (.a(c[242]), .b(s[252]), .c_in(c[243]), .s(s[678]), .c_out(c[678]));
    fullAdder fa635 (.a(s[253]), .b(c[244]), .c_in(s[254]), .s(s[679]), .c_out(c[679]));
    fullAdder fa636 (.a(c[245]), .b(s[255]), .c_in(c[246]), .s(s[680]), .c_out(c[680]));
    fullAdder fa637 (.a(s[256]), .b(c[247]), .c_in(s[257]), .s(s[681]), .c_out(c[681]));
    fullAdder fa638 (.a(c[248]), .b(s[258]), .c_in(c[249]), .s(s[682]), .c_out(c[682]));
    fullAdder fa639 (.a(s[259]), .b(c[250]), .c_in(s[260]), .s(s[683]), .c_out(c[683]));
    fullAdder fa640 (.a(c[251]), .b(s[261]), .c_in(c[252]), .s(s[684]), .c_out(c[684]));
    fullAdder fa641 (.a(s[262]), .b(c[253]), .c_in(s[263]), .s(s[685]), .c_out(c[685]));
    fullAdder fa642 (.a(c[254]), .b(s[264]), .c_in(c[255]), .s(s[686]), .c_out(c[686]));
    fullAdder fa643 (.a(s[265]), .b(c[256]), .c_in(s[266]), .s(s[687]), .c_out(c[687]));
    fullAdder fa644 (.a(c[257]), .b(s[267]), .c_in(c[258]), .s(s[688]), .c_out(c[688]));
    fullAdder fa645 (.a(s[268]), .b(c[259]), .c_in(s[269]), .s(s[689]), .c_out(c[689]));
    fullAdder fa646 (.a(c[260]), .b(s[270]), .c_in(c[261]), .s(s[690]), .c_out(c[690]));
    fullAdder fa647 (.a(s[271]), .b(c[262]), .c_in(s[272]), .s(s[691]), .c_out(c[691]));
    fullAdder fa648 (.a(c[263]), .b(s[273]), .c_in(c[264]), .s(s[692]), .c_out(c[692]));
    fullAdder fa649 (.a(s[274]), .b(c[265]), .c_in(s[275]), .s(s[693]), .c_out(c[693]));
    fullAdder fa650 (.a(c[266]), .b(s[276]), .c_in(c[267]), .s(s[694]), .c_out(c[694]));
    fullAdder fa651 (.a(s[277]), .b(c[268]), .c_in(s[278]), .s(s[695]), .c_out(c[695]));
    fullAdder fa652 (.a(c[269]), .b(s[279]), .c_in(c[270]), .s(s[696]), .c_out(c[696]));
    fullAdder fa653 (.a(s[280]), .b(c[271]), .c_in(s[281]), .s(s[697]), .c_out(c[697]));
    fullAdder fa654 (.a(c[272]), .b(s[282]), .c_in(c[273]), .s(s[698]), .c_out(c[698]));
    fullAdder fa655 (.a(s[283]), .b(c[274]), .c_in(s[284]), .s(s[699]), .c_out(c[699]));
    fullAdder fa656 (.a(c[275]), .b(s[285]), .c_in(c[276]), .s(s[700]), .c_out(c[700]));
    fullAdder fa657 (.a(s[286]), .b(c[277]), .c_in(s[287]), .s(s[701]), .c_out(c[701]));
    fullAdder fa658 (.a(c[278]), .b(s[288]), .c_in(c[279]), .s(s[702]), .c_out(c[702]));
    fullAdder fa659 (.a(s[289]), .b(c[280]), .c_in(s[290]), .s(s[703]), .c_out(c[703]));
    fullAdder fa660 (.a(c[281]), .b(s[291]), .c_in(c[282]), .s(s[704]), .c_out(c[704]));
    fullAdder fa661 (.a(s[292]), .b(c[283]), .c_in(s[293]), .s(s[705]), .c_out(c[705]));
    fullAdder fa662 (.a(c[284]), .b(s[294]), .c_in(c[285]), .s(s[706]), .c_out(c[706]));
    fullAdder fa663 (.a(s[295]), .b(c[286]), .c_in(s[296]), .s(s[707]), .c_out(c[707]));
    fullAdder fa664 (.a(c[287]), .b(s[297]), .c_in(c[288]), .s(s[708]), .c_out(c[708]));
    fullAdder fa665 (.a(s[298]), .b(c[289]), .c_in(s[299]), .s(s[709]), .c_out(c[709]));
    fullAdder fa666 (.a(c[290]), .b(s[300]), .c_in(c[291]), .s(s[710]), .c_out(c[710]));
    fullAdder fa667 (.a(s[301]), .b(c[292]), .c_in(s[302]), .s(s[711]), .c_out(c[711]));
    fullAdder fa668 (.a(c[293]), .b(p[26][06]), .c_in(c[294]), .s(s[712]), .c_out(c[712]));
    fullAdder fa669 (.a(s[303]), .b(c[295]), .c_in(s[304]), .s(s[713]), .c_out(c[713]));
    fullAdder fa670 (.a(c[296]), .b(s[305]), .c_in(c[297]), .s(s[714]), .c_out(c[714]));
    fullAdder fa671 (.a(s[306]), .b(c[298]), .c_in(s[307]), .s(s[715]), .c_out(c[715]));
    fullAdder fa672 (.a(c[299]), .b(s[308]), .c_in(c[300]), .s(s[716]), .c_out(c[716]));
    fullAdder fa673 (.a(s[309]), .b(c[301]), .c_in(s[310]), .s(s[717]), .c_out(c[717]));
    halfAdder ha46 (.a(c[302]), .b(p[26][07]), .s(s[718]), .c_out(c[718]));
    fullAdder fa674 (.a(s[311]), .b(c[303]), .c_in(s[312]), .s(s[719]), .c_out(c[719]));
    fullAdder fa675 (.a(c[304]), .b(s[313]), .c_in(c[305]), .s(s[720]), .c_out(c[720]));
    fullAdder fa676 (.a(s[314]), .b(c[306]), .c_in(s[315]), .s(s[721]), .c_out(c[721]));
    fullAdder fa677 (.a(c[307]), .b(s[316]), .c_in(c[308]), .s(s[722]), .c_out(c[722]));
    fullAdder fa678 (.a(s[317]), .b(c[309]), .c_in(s[318]), .s(s[723]), .c_out(c[723]));
    fullAdder fa679 (.a(s[319]), .b(c[311]), .c_in(s[320]), .s(s[724]), .c_out(c[724]));
    fullAdder fa680 (.a(c[312]), .b(s[321]), .c_in(c[313]), .s(s[725]), .c_out(c[725]));
    fullAdder fa681 (.a(s[322]), .b(c[314]), .c_in(s[323]), .s(s[726]), .c_out(c[726]));
    fullAdder fa682 (.a(c[315]), .b(s[324]), .c_in(c[316]), .s(s[727]), .c_out(c[727]));
    fullAdder fa683 (.a(s[325]), .b(c[317]), .c_in(s[326]), .s(s[728]), .c_out(c[728]));
    fullAdder fa684 (.a(s[327]), .b(c[319]), .c_in(s[328]), .s(s[729]), .c_out(c[729]));
    fullAdder fa685 (.a(c[320]), .b(s[329]), .c_in(c[321]), .s(s[730]), .c_out(c[730]));
    fullAdder fa686 (.a(s[330]), .b(c[322]), .c_in(s[331]), .s(s[731]), .c_out(c[731]));
    fullAdder fa687 (.a(c[323]), .b(s[332]), .c_in(c[324]), .s(s[732]), .c_out(c[732]));
    fullAdder fa688 (.a(s[333]), .b(c[325]), .c_in(s[334]), .s(s[733]), .c_out(c[733]));
    fullAdder fa689 (.a(s[335]), .b(c[327]), .c_in(s[336]), .s(s[734]), .c_out(c[734]));
    fullAdder fa690 (.a(c[328]), .b(s[337]), .c_in(c[329]), .s(s[735]), .c_out(c[735]));
    fullAdder fa691 (.a(s[338]), .b(c[330]), .c_in(s[339]), .s(s[736]), .c_out(c[736]));
    fullAdder fa692 (.a(c[331]), .b(s[340]), .c_in(c[332]), .s(s[737]), .c_out(c[737]));
    fullAdder fa693 (.a(s[341]), .b(c[333]), .c_in(s[342]), .s(s[738]), .c_out(c[738]));
    fullAdder fa694 (.a(s[343]), .b(c[335]), .c_in(s[344]), .s(s[739]), .c_out(c[739]));
    fullAdder fa695 (.a(c[336]), .b(s[345]), .c_in(c[337]), .s(s[740]), .c_out(c[740]));
    fullAdder fa696 (.a(s[346]), .b(c[338]), .c_in(s[347]), .s(s[741]), .c_out(c[741]));
    fullAdder fa697 (.a(c[339]), .b(s[348]), .c_in(c[340]), .s(s[742]), .c_out(c[742]));
    fullAdder fa698 (.a(s[349]), .b(c[341]), .c_in(p[26][12]), .s(s[743]), .c_out(c[743]));
    fullAdder fa699 (.a(s[350]), .b(c[343]), .c_in(s[351]), .s(s[744]), .c_out(c[744]));
    fullAdder fa700 (.a(c[344]), .b(s[352]), .c_in(c[345]), .s(s[745]), .c_out(c[745]));
    fullAdder fa701 (.a(s[353]), .b(c[346]), .c_in(s[354]), .s(s[746]), .c_out(c[746]));
    fullAdder fa702 (.a(c[347]), .b(s[355]), .c_in(c[348]), .s(s[747]), .c_out(c[747]));
    fullAdder fa703 (.a(s[356]), .b(c[349]), .c_in(p[26][13]), .s(s[748]), .c_out(c[748]));
    fullAdder fa704 (.a(s[357]), .b(c[350]), .c_in(s[358]), .s(s[749]), .c_out(c[749]));
    fullAdder fa705 (.a(c[351]), .b(s[359]), .c_in(c[352]), .s(s[750]), .c_out(c[750]));
    fullAdder fa706 (.a(s[360]), .b(c[353]), .c_in(s[361]), .s(s[751]), .c_out(c[751]));
    fullAdder fa707 (.a(c[354]), .b(s[362]), .c_in(c[355]), .s(s[752]), .c_out(c[752]));
    halfAdder ha47 (.a(s[363]), .b(c[356]), .s(s[753]), .c_out(c[753]));
    fullAdder fa708 (.a(s[364]), .b(c[357]), .c_in(s[365]), .s(s[754]), .c_out(c[754]));
    fullAdder fa709 (.a(c[358]), .b(s[366]), .c_in(c[359]), .s(s[755]), .c_out(c[755]));
    fullAdder fa710 (.a(s[367]), .b(c[360]), .c_in(s[368]), .s(s[756]), .c_out(c[756]));
    fullAdder fa711 (.a(c[361]), .b(s[369]), .c_in(c[362]), .s(s[757]), .c_out(c[757]));
    halfAdder ha48 (.a(s[370]), .b(c[363]), .s(s[758]), .c_out(c[758]));
    fullAdder fa712 (.a(s[371]), .b(c[364]), .c_in(s[372]), .s(s[759]), .c_out(c[759]));
    fullAdder fa713 (.a(c[365]), .b(s[373]), .c_in(c[366]), .s(s[760]), .c_out(c[760]));
    fullAdder fa714 (.a(s[374]), .b(c[367]), .c_in(s[375]), .s(s[761]), .c_out(c[761]));
    fullAdder fa715 (.a(c[368]), .b(s[376]), .c_in(c[369]), .s(s[762]), .c_out(c[762]));
    halfAdder ha49 (.a(s[377]), .b(c[370]), .s(s[763]), .c_out(c[763]));
    fullAdder fa716 (.a(s[378]), .b(c[371]), .c_in(s[379]), .s(s[764]), .c_out(c[764]));
    fullAdder fa717 (.a(c[372]), .b(s[380]), .c_in(c[373]), .s(s[765]), .c_out(c[765]));
    fullAdder fa718 (.a(s[381]), .b(c[374]), .c_in(s[382]), .s(s[766]), .c_out(c[766]));
    fullAdder fa719 (.a(c[375]), .b(s[383]), .c_in(c[376]), .s(s[767]), .c_out(c[767]));
    halfAdder ha50 (.a(s[384]), .b(c[377]), .s(s[768]), .c_out(c[768]));
    fullAdder fa720 (.a(s[385]), .b(c[378]), .c_in(s[386]), .s(s[769]), .c_out(c[769]));
    fullAdder fa721 (.a(c[379]), .b(s[387]), .c_in(c[380]), .s(s[770]), .c_out(c[770]));
    fullAdder fa722 (.a(s[388]), .b(c[381]), .c_in(s[389]), .s(s[771]), .c_out(c[771]));
    fullAdder fa723 (.a(c[382]), .b(s[390]), .c_in(c[383]), .s(s[772]), .c_out(c[772]));
    halfAdder ha51 (.a(p[26][18]), .b(c[384]), .s(s[773]), .c_out(c[773]));
    fullAdder fa724 (.a(s[391]), .b(c[385]), .c_in(s[392]), .s(s[774]), .c_out(c[774]));
    fullAdder fa725 (.a(c[386]), .b(s[393]), .c_in(c[387]), .s(s[775]), .c_out(c[775]));
    fullAdder fa726 (.a(s[394]), .b(c[388]), .c_in(s[395]), .s(s[776]), .c_out(c[776]));
    fullAdder fa727 (.a(c[389]), .b(s[396]), .c_in(c[390]), .s(s[777]), .c_out(c[777]));
    fullAdder fa728 (.a(s[397]), .b(c[391]), .c_in(s[398]), .s(s[778]), .c_out(c[778]));
    fullAdder fa729 (.a(c[392]), .b(s[399]), .c_in(c[393]), .s(s[779]), .c_out(c[779]));
    fullAdder fa730 (.a(s[400]), .b(c[394]), .c_in(s[401]), .s(s[780]), .c_out(c[780]));
    fullAdder fa731 (.a(c[395]), .b(s[402]), .c_in(c[396]), .s(s[781]), .c_out(c[781]));
    fullAdder fa732 (.a(s[403]), .b(c[397]), .c_in(s[404]), .s(s[782]), .c_out(c[782]));
    fullAdder fa733 (.a(c[398]), .b(s[405]), .c_in(c[399]), .s(s[783]), .c_out(c[783]));
    fullAdder fa734 (.a(s[406]), .b(c[400]), .c_in(s[407]), .s(s[784]), .c_out(c[784]));
    fullAdder fa735 (.a(c[401]), .b(s[408]), .c_in(c[402]), .s(s[785]), .c_out(c[785]));
    fullAdder fa736 (.a(s[409]), .b(c[403]), .c_in(s[410]), .s(s[786]), .c_out(c[786]));
    fullAdder fa737 (.a(c[404]), .b(s[411]), .c_in(c[405]), .s(s[787]), .c_out(c[787]));
    fullAdder fa738 (.a(s[412]), .b(c[406]), .c_in(s[413]), .s(s[788]), .c_out(c[788]));
    fullAdder fa739 (.a(c[407]), .b(s[414]), .c_in(c[408]), .s(s[789]), .c_out(c[789]));
    fullAdder fa740 (.a(s[415]), .b(c[409]), .c_in(s[416]), .s(s[790]), .c_out(c[790]));
    fullAdder fa741 (.a(c[410]), .b(s[417]), .c_in(c[411]), .s(s[791]), .c_out(c[791]));
    fullAdder fa742 (.a(s[418]), .b(c[412]), .c_in(s[419]), .s(s[792]), .c_out(c[792]));
    fullAdder fa743 (.a(c[413]), .b(s[420]), .c_in(c[414]), .s(s[793]), .c_out(c[793]));
    fullAdder fa744 (.a(s[421]), .b(c[415]), .c_in(s[422]), .s(s[794]), .c_out(c[794]));
    fullAdder fa745 (.a(c[416]), .b(s[423]), .c_in(c[417]), .s(s[795]), .c_out(c[795]));
    fullAdder fa746 (.a(s[424]), .b(c[418]), .c_in(s[425]), .s(s[796]), .c_out(c[796]));
    fullAdder fa747 (.a(c[419]), .b(p[26][24]), .c_in(c[420]), .s(s[797]), .c_out(c[797]));
    fullAdder fa748 (.a(s[426]), .b(c[421]), .c_in(s[427]), .s(s[798]), .c_out(c[798]));
    fullAdder fa749 (.a(c[422]), .b(s[428]), .c_in(c[423]), .s(s[799]), .c_out(c[799]));
    fullAdder fa750 (.a(s[429]), .b(c[424]), .c_in(s[430]), .s(s[800]), .c_out(c[800]));
    halfAdder ha52 (.a(c[425]), .b(p[26][25]), .s(s[801]), .c_out(c[801]));
    fullAdder fa751 (.a(s[431]), .b(c[426]), .c_in(s[432]), .s(s[802]), .c_out(c[802]));
    fullAdder fa752 (.a(c[427]), .b(s[433]), .c_in(c[428]), .s(s[803]), .c_out(c[803]));
    fullAdder fa753 (.a(s[434]), .b(c[429]), .c_in(s[435]), .s(s[804]), .c_out(c[804]));
    fullAdder fa754 (.a(s[436]), .b(c[431]), .c_in(s[437]), .s(s[805]), .c_out(c[805]));
    fullAdder fa755 (.a(c[432]), .b(s[438]), .c_in(c[433]), .s(s[806]), .c_out(c[806]));
    fullAdder fa756 (.a(s[439]), .b(c[434]), .c_in(s[440]), .s(s[807]), .c_out(c[807]));
    fullAdder fa757 (.a(s[441]), .b(c[436]), .c_in(s[442]), .s(s[808]), .c_out(c[808]));
    fullAdder fa758 (.a(c[437]), .b(s[443]), .c_in(c[438]), .s(s[809]), .c_out(c[809]));
    fullAdder fa759 (.a(s[444]), .b(c[439]), .c_in(s[445]), .s(s[810]), .c_out(c[810]));
    fullAdder fa760 (.a(s[446]), .b(c[441]), .c_in(s[447]), .s(s[811]), .c_out(c[811]));
    fullAdder fa761 (.a(c[442]), .b(s[448]), .c_in(c[443]), .s(s[812]), .c_out(c[812]));
    fullAdder fa762 (.a(s[449]), .b(c[444]), .c_in(s[450]), .s(s[813]), .c_out(c[813]));
    fullAdder fa763 (.a(s[451]), .b(c[446]), .c_in(s[452]), .s(s[814]), .c_out(c[814]));
    fullAdder fa764 (.a(c[447]), .b(s[453]), .c_in(c[448]), .s(s[815]), .c_out(c[815]));
    fullAdder fa765 (.a(s[454]), .b(c[449]), .c_in(p[26][30]), .s(s[816]), .c_out(c[816]));
    fullAdder fa766 (.a(s[455]), .b(c[451]), .c_in(s[456]), .s(s[817]), .c_out(c[817]));
    fullAdder fa767 (.a(c[452]), .b(s[457]), .c_in(c[453]), .s(s[818]), .c_out(c[818]));
    fullAdder fa768 (.a(s[458]), .b(c[454]), .c_in(p[26][31]), .s(s[819]), .c_out(c[819]));
    fullAdder fa769 (.a(s[459]), .b(c[455]), .c_in(s[460]), .s(s[820]), .c_out(c[820]));
    fullAdder fa770 (.a(c[456]), .b(s[461]), .c_in(c[457]), .s(s[821]), .c_out(c[821]));
    fullAdder fa771 (.a(s[462]), .b(c[458]), .c_in(p[26][32]), .s(s[822]), .c_out(c[822]));
    fullAdder fa772 (.a(s[463]), .b(c[459]), .c_in(s[464]), .s(s[823]), .c_out(c[823]));
    fullAdder fa773 (.a(c[460]), .b(s[465]), .c_in(c[461]), .s(s[824]), .c_out(c[824]));
    halfAdder ha53 (.a(s[466]), .b(c[462]), .s(s[825]), .c_out(c[825]));
    fullAdder fa774 (.a(s[467]), .b(c[463]), .c_in(s[468]), .s(s[826]), .c_out(c[826]));
    fullAdder fa775 (.a(c[464]), .b(s[469]), .c_in(c[465]), .s(s[827]), .c_out(c[827]));
    halfAdder ha54 (.a(s[470]), .b(c[466]), .s(s[828]), .c_out(c[828]));
    fullAdder fa776 (.a(s[471]), .b(c[467]), .c_in(s[472]), .s(s[829]), .c_out(c[829]));
    fullAdder fa777 (.a(c[468]), .b(s[473]), .c_in(c[469]), .s(s[830]), .c_out(c[830]));
    halfAdder ha55 (.a(s[474]), .b(c[470]), .s(s[831]), .c_out(c[831]));
    fullAdder fa778 (.a(s[475]), .b(c[471]), .c_in(s[476]), .s(s[832]), .c_out(c[832]));
    fullAdder fa779 (.a(c[472]), .b(s[477]), .c_in(c[473]), .s(s[833]), .c_out(c[833]));
    halfAdder ha56 (.a(p[26][36]), .b(c[474]), .s(s[834]), .c_out(c[834]));
    fullAdder fa780 (.a(s[478]), .b(c[475]), .c_in(s[479]), .s(s[835]), .c_out(c[835]));
    fullAdder fa781 (.a(c[476]), .b(s[480]), .c_in(c[477]), .s(s[836]), .c_out(c[836]));
    fullAdder fa782 (.a(s[481]), .b(c[478]), .c_in(s[482]), .s(s[837]), .c_out(c[837]));
    fullAdder fa783 (.a(c[479]), .b(s[483]), .c_in(c[480]), .s(s[838]), .c_out(c[838]));
    fullAdder fa784 (.a(s[484]), .b(c[481]), .c_in(s[485]), .s(s[839]), .c_out(c[839]));
    fullAdder fa785 (.a(c[482]), .b(s[486]), .c_in(c[483]), .s(s[840]), .c_out(c[840]));
    fullAdder fa786 (.a(s[487]), .b(c[484]), .c_in(s[488]), .s(s[841]), .c_out(c[841]));
    fullAdder fa787 (.a(c[485]), .b(s[489]), .c_in(c[486]), .s(s[842]), .c_out(c[842]));
    fullAdder fa788 (.a(s[490]), .b(c[487]), .c_in(s[491]), .s(s[843]), .c_out(c[843]));
    fullAdder fa789 (.a(c[488]), .b(s[492]), .c_in(c[489]), .s(s[844]), .c_out(c[844]));
    fullAdder fa790 (.a(s[493]), .b(c[490]), .c_in(s[494]), .s(s[845]), .c_out(c[845]));
    fullAdder fa791 (.a(c[491]), .b(p[26][42]), .c_in(c[492]), .s(s[846]), .c_out(c[846]));
    fullAdder fa792 (.a(s[495]), .b(c[493]), .c_in(s[496]), .s(s[847]), .c_out(c[847]));
    halfAdder ha57 (.a(c[494]), .b(p[26][43]), .s(s[848]), .c_out(c[848]));
    fullAdder fa793 (.a(s[497]), .b(c[495]), .c_in(s[498]), .s(s[849]), .c_out(c[849]));
    fullAdder fa794 (.a(s[499]), .b(c[497]), .c_in(s[500]), .s(s[850]), .c_out(c[850]));
    fullAdder fa795 (.a(s[501]), .b(c[499]), .c_in(s[502]), .s(s[851]), .c_out(c[851]));
    fullAdder fa796 (.a(s[503]), .b(c[501]), .c_in(s[504]), .s(s[852]), .c_out(c[852]));
    fullAdder fa797 (.a(s[505]), .b(c[503]), .c_in(p[26][48]), .s(s[853]), .c_out(c[853]));
    fullAdder fa798 (.a(s[506]), .b(c[505]), .c_in(p[26][49]), .s(s[854]), .c_out(c[854]));
    fullAdder fa799 (.a(~comp[25]), .b(c[508]), .c_in(p[26][52]), .s(s[855]), .c_out(c[855]));
    // Stage 3 Reduction
    fullAdder fa800 (.a(s[1]), .b(c[509]), .c_in(comp[2]), .s(s[856]), .c_out(c[856]));
    fullAdder fa801 (.a(s[511]), .b(c[510]), .c_in(c[4]), .s(s[857]), .c_out(c[857]));
    fullAdder fa802 (.a(s[513]), .b(c[512]), .c_in(c[7]), .s(s[858]), .c_out(c[858]));
    fullAdder fa803 (.a(s[514]), .b(c[513]), .c_in(s[515]), .s(s[859]), .c_out(c[859]));
    fullAdder fa804 (.a(s[516]), .b(c[514]), .c_in(c[11]), .s(s[860]), .c_out(c[860]));
    fullAdder fa805 (.a(s[517]), .b(c[516]), .c_in(s[518]), .s(s[861]), .c_out(c[861]));
    fullAdder fa806 (.a(s[519]), .b(c[517]), .c_in(s[520]), .s(s[862]), .c_out(c[862]));
    fullAdder fa807 (.a(s[521]), .b(c[519]), .c_in(s[522]), .s(s[863]), .c_out(c[863]));
    fullAdder fa808 (.a(s[523]), .b(c[521]), .c_in(s[524]), .s(s[864]), .c_out(c[864]));
    fullAdder fa809 (.a(s[525]), .b(c[523]), .c_in(s[526]), .s(s[865]), .c_out(c[865]));
    halfAdder ha58 (.a(c[524]), .b(mode == 2'b01 ? 1'b0 : comp[8]), .s(s[866]), .c_out(c[866]));
    fullAdder fa810 (.a(s[527]), .b(c[525]), .c_in(s[528]), .s(s[867]), .c_out(c[867]));
    fullAdder fa811 (.a(s[529]), .b(c[527]), .c_in(s[530]), .s(s[868]), .c_out(c[868]));
    halfAdder ha59 (.a(c[528]), .b(s[34]), .s(s[869]), .c_out(c[869]));
    fullAdder fa812 (.a(s[531]), .b(c[529]), .c_in(s[532]), .s(s[870]), .c_out(c[870]));
    halfAdder ha60 (.a(c[530]), .b(s[533]), .s(s[871]), .c_out(c[871]));
    fullAdder fa813 (.a(s[534]), .b(c[531]), .c_in(s[535]), .s(s[872]), .c_out(c[872]));
    fullAdder fa814 (.a(c[532]), .b(s[41]), .c_in(c[533]), .s(s[873]), .c_out(c[873]));
    fullAdder fa815 (.a(s[536]), .b(c[534]), .c_in(s[537]), .s(s[874]), .c_out(c[874]));
    halfAdder ha61 (.a(c[535]), .b(s[538]), .s(s[875]), .c_out(c[875]));
    fullAdder fa816 (.a(s[539]), .b(c[536]), .c_in(s[540]), .s(s[876]), .c_out(c[876]));
    fullAdder fa817 (.a(c[537]), .b(s[541]), .c_in(c[538]), .s(s[877]), .c_out(c[877]));
    fullAdder fa818 (.a(s[542]), .b(c[539]), .c_in(s[543]), .s(s[878]), .c_out(c[878]));
    fullAdder fa819 (.a(c[540]), .b(s[544]), .c_in(c[541]), .s(s[879]), .c_out(c[879]));
    fullAdder fa820 (.a(s[545]), .b(c[542]), .c_in(s[546]), .s(s[880]), .c_out(c[880]));
    fullAdder fa821 (.a(c[543]), .b(s[547]), .c_in(c[544]), .s(s[881]), .c_out(c[881]));
    fullAdder fa822 (.a(s[548]), .b(c[545]), .c_in(s[549]), .s(s[882]), .c_out(c[882]));
    fullAdder fa823 (.a(c[546]), .b(s[550]), .c_in(c[547]), .s(s[883]), .c_out(c[883]));
    fullAdder fa824 (.a(s[551]), .b(c[548]), .c_in(s[552]), .s(s[884]), .c_out(c[884]));
    fullAdder fa825 (.a(c[549]), .b(s[553]), .c_in(c[550]), .s(s[885]), .c_out(c[885]));
    fullAdder fa826 (.a(s[554]), .b(c[551]), .c_in(s[555]), .s(s[886]), .c_out(c[886]));
    fullAdder fa827 (.a(c[552]), .b(s[556]), .c_in(c[553]), .s(s[887]), .c_out(c[887]));
    fullAdder fa828 (.a(s[557]), .b(c[554]), .c_in(s[558]), .s(s[888]), .c_out(c[888]));
    fullAdder fa829 (.a(c[555]), .b(s[559]), .c_in(c[556]), .s(s[889]), .c_out(c[889]));
    fullAdder fa830 (.a(s[561]), .b(c[557]), .c_in(s[562]), .s(s[890]), .c_out(c[890]));
    fullAdder fa831 (.a(c[558]), .b(s[563]), .c_in(c[559]), .s(s[891]), .c_out(c[891]));
    halfAdder ha62 (.a(c[77]), .b(c[560]), .s(s[892]), .c_out(c[892]));
    fullAdder fa832 (.a(s[564]), .b(c[561]), .c_in(s[565]), .s(s[893]), .c_out(c[893]));
    fullAdder fa833 (.a(c[562]), .b(s[566]), .c_in(c[563]), .s(s[894]), .c_out(c[894]));
    fullAdder fa834 (.a(s[568]), .b(c[564]), .c_in(s[569]), .s(s[895]), .c_out(c[895]));
    fullAdder fa835 (.a(c[565]), .b(s[570]), .c_in(c[566]), .s(s[896]), .c_out(c[896]));
    halfAdder ha63 (.a(s[571]), .b(c[567]), .s(s[897]), .c_out(c[897]));
    fullAdder fa836 (.a(s[572]), .b(c[568]), .c_in(s[573]), .s(s[898]), .c_out(c[898]));
    fullAdder fa837 (.a(c[569]), .b(s[574]), .c_in(c[570]), .s(s[899]), .c_out(c[899]));
    halfAdder ha64 (.a(s[575]), .b(c[571]), .s(s[900]), .c_out(c[900]));
    fullAdder fa838 (.a(s[576]), .b(c[572]), .c_in(s[577]), .s(s[901]), .c_out(c[901]));
    fullAdder fa839 (.a(c[573]), .b(s[578]), .c_in(c[574]), .s(s[902]), .c_out(c[902]));
    halfAdder ha65 (.a(s[579]), .b(c[575]), .s(s[903]), .c_out(c[903]));
    fullAdder fa840 (.a(s[580]), .b(c[576]), .c_in(s[581]), .s(s[904]), .c_out(c[904]));
    fullAdder fa841 (.a(c[577]), .b(s[582]), .c_in(c[578]), .s(s[905]), .c_out(c[905]));
    fullAdder fa842 (.a(s[583]), .b(c[579]), .c_in(mode == 2'b11 ? comp[17] : 1'b0), .s(s[906]), .c_out(c[906]));
    fullAdder fa843 (.a(s[584]), .b(c[580]), .c_in(s[585]), .s(s[907]), .c_out(c[907]));
    fullAdder fa844 (.a(c[581]), .b(s[586]), .c_in(c[582]), .s(s[908]), .c_out(c[908]));
    halfAdder ha66 (.a(s[587]), .b(c[583]), .s(s[909]), .c_out(c[909]));
    fullAdder fa845 (.a(s[588]), .b(c[584]), .c_in(s[589]), .s(s[910]), .c_out(c[910]));
    fullAdder fa846 (.a(c[585]), .b(s[590]), .c_in(c[586]), .s(s[911]), .c_out(c[911]));
    fullAdder fa847 (.a(s[591]), .b(c[587]), .c_in(s[124]), .s(s[912]), .c_out(c[912]));
    fullAdder fa848 (.a(s[592]), .b(c[588]), .c_in(s[593]), .s(s[913]), .c_out(c[913]));
    fullAdder fa849 (.a(c[589]), .b(s[594]), .c_in(c[590]), .s(s[914]), .c_out(c[914]));
    fullAdder fa850 (.a(s[595]), .b(c[591]), .c_in(s[596]), .s(s[915]), .c_out(c[915]));
    fullAdder fa851 (.a(s[597]), .b(c[592]), .c_in(s[598]), .s(s[916]), .c_out(c[916]));
    fullAdder fa852 (.a(c[593]), .b(s[599]), .c_in(c[594]), .s(s[917]), .c_out(c[917]));
    fullAdder fa853 (.a(s[600]), .b(c[595]), .c_in(s[137]), .s(s[918]), .c_out(c[918]));
    fullAdder fa854 (.a(s[601]), .b(c[597]), .c_in(s[602]), .s(s[919]), .c_out(c[919]));
    fullAdder fa855 (.a(c[598]), .b(s[603]), .c_in(c[599]), .s(s[920]), .c_out(c[920]));
    fullAdder fa856 (.a(s[604]), .b(c[600]), .c_in(s[605]), .s(s[921]), .c_out(c[921]));
    fullAdder fa857 (.a(s[606]), .b(c[601]), .c_in(s[607]), .s(s[922]), .c_out(c[922]));
    fullAdder fa858 (.a(c[602]), .b(s[608]), .c_in(c[603]), .s(s[923]), .c_out(c[923]));
    fullAdder fa859 (.a(s[609]), .b(c[604]), .c_in(s[610]), .s(s[924]), .c_out(c[924]));
    fullAdder fa860 (.a(s[611]), .b(c[606]), .c_in(s[612]), .s(s[925]), .c_out(c[925]));
    fullAdder fa861 (.a(c[607]), .b(s[613]), .c_in(c[608]), .s(s[926]), .c_out(c[926]));
    fullAdder fa862 (.a(s[614]), .b(c[609]), .c_in(s[615]), .s(s[927]), .c_out(c[927]));
    fullAdder fa863 (.a(s[616]), .b(c[611]), .c_in(s[617]), .s(s[928]), .c_out(c[928]));
    fullAdder fa864 (.a(c[612]), .b(s[618]), .c_in(c[613]), .s(s[929]), .c_out(c[929]));
    fullAdder fa865 (.a(s[619]), .b(c[614]), .c_in(s[620]), .s(s[930]), .c_out(c[930]));
    fullAdder fa866 (.a(s[621]), .b(c[616]), .c_in(s[622]), .s(s[931]), .c_out(c[931]));
    fullAdder fa867 (.a(c[617]), .b(s[623]), .c_in(c[618]), .s(s[932]), .c_out(c[932]));
    fullAdder fa868 (.a(s[624]), .b(c[619]), .c_in(s[625]), .s(s[933]), .c_out(c[933]));
    halfAdder ha67 (.a(c[620]), .b(c[166]), .s(s[934]), .c_out(c[934]));
    fullAdder fa869 (.a(s[626]), .b(c[621]), .c_in(s[627]), .s(s[935]), .c_out(c[935]));
    fullAdder fa870 (.a(c[622]), .b(s[628]), .c_in(c[623]), .s(s[936]), .c_out(c[936]));
    fullAdder fa871 (.a(s[629]), .b(c[624]), .c_in(s[630]), .s(s[937]), .c_out(c[937]));
    fullAdder fa872 (.a(s[631]), .b(c[626]), .c_in(s[632]), .s(s[938]), .c_out(c[938]));
    fullAdder fa873 (.a(c[627]), .b(s[633]), .c_in(c[628]), .s(s[939]), .c_out(c[939]));
    fullAdder fa874 (.a(s[634]), .b(c[629]), .c_in(s[635]), .s(s[940]), .c_out(c[940]));
    halfAdder ha68 (.a(c[630]), .b(c[181]), .s(s[941]), .c_out(c[941]));
    fullAdder fa875 (.a(s[636]), .b(c[631]), .c_in(s[637]), .s(s[942]), .c_out(c[942]));
    fullAdder fa876 (.a(c[632]), .b(s[638]), .c_in(c[633]), .s(s[943]), .c_out(c[943]));
    fullAdder fa877 (.a(s[639]), .b(c[634]), .c_in(s[640]), .s(s[944]), .c_out(c[944]));
    halfAdder ha69 (.a(c[635]), .b(s[641]), .s(s[945]), .c_out(c[945]));
    fullAdder fa878 (.a(s[642]), .b(c[636]), .c_in(s[643]), .s(s[946]), .c_out(c[946]));
    fullAdder fa879 (.a(c[637]), .b(s[644]), .c_in(c[638]), .s(s[947]), .c_out(c[947]));
    fullAdder fa880 (.a(s[645]), .b(c[639]), .c_in(s[646]), .s(s[948]), .c_out(c[948]));
    fullAdder fa881 (.a(c[640]), .b(c[197]), .c_in(c[641]), .s(s[949]), .c_out(c[949]));
    fullAdder fa882 (.a(s[647]), .b(c[642]), .c_in(s[648]), .s(s[950]), .c_out(c[950]));
    fullAdder fa883 (.a(c[643]), .b(s[649]), .c_in(c[644]), .s(s[951]), .c_out(c[951]));
    fullAdder fa884 (.a(s[650]), .b(c[645]), .c_in(s[651]), .s(s[952]), .c_out(c[952]));
    halfAdder ha70 (.a(c[646]), .b(s[652]), .s(s[953]), .c_out(c[953]));
    fullAdder fa885 (.a(s[653]), .b(c[647]), .c_in(s[654]), .s(s[954]), .c_out(c[954]));
    fullAdder fa886 (.a(c[648]), .b(s[655]), .c_in(c[649]), .s(s[955]), .c_out(c[955]));
    fullAdder fa887 (.a(s[656]), .b(c[650]), .c_in(s[657]), .s(s[956]), .c_out(c[956]));
    fullAdder fa888 (.a(c[651]), .b(s[658]), .c_in(c[652]), .s(s[957]), .c_out(c[957]));
    fullAdder fa889 (.a(s[659]), .b(c[653]), .c_in(s[660]), .s(s[958]), .c_out(c[958]));
    fullAdder fa890 (.a(c[654]), .b(s[661]), .c_in(c[655]), .s(s[959]), .c_out(c[959]));
    fullAdder fa891 (.a(s[662]), .b(c[656]), .c_in(s[663]), .s(s[960]), .c_out(c[960]));
    fullAdder fa892 (.a(c[657]), .b(s[664]), .c_in(c[658]), .s(s[961]), .c_out(c[961]));
    fullAdder fa893 (.a(s[665]), .b(c[659]), .c_in(s[666]), .s(s[962]), .c_out(c[962]));
    fullAdder fa894 (.a(c[660]), .b(s[667]), .c_in(c[661]), .s(s[963]), .c_out(c[963]));
    fullAdder fa895 (.a(s[668]), .b(c[662]), .c_in(s[669]), .s(s[964]), .c_out(c[964]));
    fullAdder fa896 (.a(c[663]), .b(s[670]), .c_in(c[664]), .s(s[965]), .c_out(c[965]));
    fullAdder fa897 (.a(s[671]), .b(c[665]), .c_in(s[672]), .s(s[966]), .c_out(c[966]));
    fullAdder fa898 (.a(c[666]), .b(s[673]), .c_in(c[667]), .s(s[967]), .c_out(c[967]));
    fullAdder fa899 (.a(s[674]), .b(c[668]), .c_in(s[675]), .s(s[968]), .c_out(c[968]));
    fullAdder fa900 (.a(c[669]), .b(s[676]), .c_in(c[670]), .s(s[969]), .c_out(c[969]));
    fullAdder fa901 (.a(s[677]), .b(c[671]), .c_in(s[678]), .s(s[970]), .c_out(c[970]));
    fullAdder fa902 (.a(c[672]), .b(s[679]), .c_in(c[673]), .s(s[971]), .c_out(c[971]));
    fullAdder fa903 (.a(s[680]), .b(c[674]), .c_in(s[681]), .s(s[972]), .c_out(c[972]));
    fullAdder fa904 (.a(c[675]), .b(s[682]), .c_in(c[676]), .s(s[973]), .c_out(c[973]));
    fullAdder fa905 (.a(s[683]), .b(c[677]), .c_in(s[684]), .s(s[974]), .c_out(c[974]));
    fullAdder fa906 (.a(c[678]), .b(s[685]), .c_in(c[679]), .s(s[975]), .c_out(c[975]));
    fullAdder fa907 (.a(s[686]), .b(c[680]), .c_in(s[687]), .s(s[976]), .c_out(c[976]));
    fullAdder fa908 (.a(c[681]), .b(s[688]), .c_in(c[682]), .s(s[977]), .c_out(c[977]));
    fullAdder fa909 (.a(s[689]), .b(c[683]), .c_in(s[690]), .s(s[978]), .c_out(c[978]));
    fullAdder fa910 (.a(c[684]), .b(s[691]), .c_in(c[685]), .s(s[979]), .c_out(c[979]));
    fullAdder fa911 (.a(s[692]), .b(c[686]), .c_in(s[693]), .s(s[980]), .c_out(c[980]));
    fullAdder fa912 (.a(c[687]), .b(s[694]), .c_in(c[688]), .s(s[981]), .c_out(c[981]));
    fullAdder fa913 (.a(s[695]), .b(c[689]), .c_in(s[696]), .s(s[982]), .c_out(c[982]));
    fullAdder fa914 (.a(c[690]), .b(s[697]), .c_in(c[691]), .s(s[983]), .c_out(c[983]));
    fullAdder fa915 (.a(s[698]), .b(c[692]), .c_in(s[699]), .s(s[984]), .c_out(c[984]));
    fullAdder fa916 (.a(c[693]), .b(s[700]), .c_in(c[694]), .s(s[985]), .c_out(c[985]));
    fullAdder fa917 (.a(s[701]), .b(c[695]), .c_in(s[702]), .s(s[986]), .c_out(c[986]));
    fullAdder fa918 (.a(c[696]), .b(s[703]), .c_in(c[697]), .s(s[987]), .c_out(c[987]));
    fullAdder fa919 (.a(s[704]), .b(c[698]), .c_in(s[705]), .s(s[988]), .c_out(c[988]));
    fullAdder fa920 (.a(c[699]), .b(s[706]), .c_in(c[700]), .s(s[989]), .c_out(c[989]));
    fullAdder fa921 (.a(s[707]), .b(c[701]), .c_in(s[708]), .s(s[990]), .c_out(c[990]));
    fullAdder fa922 (.a(c[702]), .b(s[709]), .c_in(c[703]), .s(s[991]), .c_out(c[991]));
    fullAdder fa923 (.a(s[710]), .b(c[704]), .c_in(s[711]), .s(s[992]), .c_out(c[992]));
    fullAdder fa924 (.a(c[705]), .b(s[712]), .c_in(c[706]), .s(s[993]), .c_out(c[993]));
    fullAdder fa925 (.a(s[713]), .b(c[707]), .c_in(s[714]), .s(s[994]), .c_out(c[994]));
    fullAdder fa926 (.a(c[708]), .b(s[715]), .c_in(c[709]), .s(s[995]), .c_out(c[995]));
    fullAdder fa927 (.a(s[716]), .b(c[710]), .c_in(s[717]), .s(s[996]), .c_out(c[996]));
    fullAdder fa928 (.a(c[711]), .b(s[718]), .c_in(c[712]), .s(s[997]), .c_out(c[997]));
    fullAdder fa929 (.a(s[719]), .b(c[713]), .c_in(s[720]), .s(s[998]), .c_out(c[998]));
    fullAdder fa930 (.a(c[714]), .b(s[721]), .c_in(c[715]), .s(s[999]), .c_out(c[999]));
    fullAdder fa931 (.a(s[722]), .b(c[716]), .c_in(s[723]), .s(s[1000]), .c_out(c[1000]));
    fullAdder fa932 (.a(c[717]), .b(c[310]), .c_in(c[718]), .s(s[1001]), .c_out(c[1001]));
    fullAdder fa933 (.a(s[724]), .b(c[719]), .c_in(s[725]), .s(s[1002]), .c_out(c[1002]));
    fullAdder fa934 (.a(c[720]), .b(s[726]), .c_in(c[721]), .s(s[1003]), .c_out(c[1003]));
    fullAdder fa935 (.a(s[727]), .b(c[722]), .c_in(s[728]), .s(s[1004]), .c_out(c[1004]));
    halfAdder ha71 (.a(c[723]), .b(c[318]), .s(s[1005]), .c_out(c[1005]));
    fullAdder fa936 (.a(s[729]), .b(c[724]), .c_in(s[730]), .s(s[1006]), .c_out(c[1006]));
    fullAdder fa937 (.a(c[725]), .b(s[731]), .c_in(c[726]), .s(s[1007]), .c_out(c[1007]));
    fullAdder fa938 (.a(s[732]), .b(c[727]), .c_in(s[733]), .s(s[1008]), .c_out(c[1008]));
    halfAdder ha72 (.a(c[728]), .b(c[326]), .s(s[1009]), .c_out(c[1009]));
    fullAdder fa939 (.a(s[734]), .b(c[729]), .c_in(s[735]), .s(s[1010]), .c_out(c[1010]));
    fullAdder fa940 (.a(c[730]), .b(s[736]), .c_in(c[731]), .s(s[1011]), .c_out(c[1011]));
    fullAdder fa941 (.a(s[737]), .b(c[732]), .c_in(s[738]), .s(s[1012]), .c_out(c[1012]));
    halfAdder ha73 (.a(c[733]), .b(c[334]), .s(s[1013]), .c_out(c[1013]));
    fullAdder fa942 (.a(s[739]), .b(c[734]), .c_in(s[740]), .s(s[1014]), .c_out(c[1014]));
    fullAdder fa943 (.a(c[735]), .b(s[741]), .c_in(c[736]), .s(s[1015]), .c_out(c[1015]));
    fullAdder fa944 (.a(s[742]), .b(c[737]), .c_in(s[743]), .s(s[1016]), .c_out(c[1016]));
    halfAdder ha74 (.a(c[738]), .b(c[342]), .s(s[1017]), .c_out(c[1017]));
    fullAdder fa945 (.a(s[744]), .b(c[739]), .c_in(s[745]), .s(s[1018]), .c_out(c[1018]));
    fullAdder fa946 (.a(c[740]), .b(s[746]), .c_in(c[741]), .s(s[1019]), .c_out(c[1019]));
    fullAdder fa947 (.a(s[747]), .b(c[742]), .c_in(s[748]), .s(s[1020]), .c_out(c[1020]));
    fullAdder fa948 (.a(s[749]), .b(c[744]), .c_in(s[750]), .s(s[1021]), .c_out(c[1021]));
    fullAdder fa949 (.a(c[745]), .b(s[751]), .c_in(c[746]), .s(s[1022]), .c_out(c[1022]));
    fullAdder fa950 (.a(s[752]), .b(c[747]), .c_in(s[753]), .s(s[1023]), .c_out(c[1023]));
    fullAdder fa951 (.a(s[754]), .b(c[749]), .c_in(s[755]), .s(s[1024]), .c_out(c[1024]));
    fullAdder fa952 (.a(c[750]), .b(s[756]), .c_in(c[751]), .s(s[1025]), .c_out(c[1025]));
    fullAdder fa953 (.a(s[757]), .b(c[752]), .c_in(s[758]), .s(s[1026]), .c_out(c[1026]));
    fullAdder fa954 (.a(s[759]), .b(c[754]), .c_in(s[760]), .s(s[1027]), .c_out(c[1027]));
    fullAdder fa955 (.a(c[755]), .b(s[761]), .c_in(c[756]), .s(s[1028]), .c_out(c[1028]));
    fullAdder fa956 (.a(s[762]), .b(c[757]), .c_in(s[763]), .s(s[1029]), .c_out(c[1029]));
    fullAdder fa957 (.a(s[764]), .b(c[759]), .c_in(s[765]), .s(s[1030]), .c_out(c[1030]));
    fullAdder fa958 (.a(c[760]), .b(s[766]), .c_in(c[761]), .s(s[1031]), .c_out(c[1031]));
    fullAdder fa959 (.a(s[767]), .b(c[762]), .c_in(s[768]), .s(s[1032]), .c_out(c[1032]));
    fullAdder fa960 (.a(s[769]), .b(c[764]), .c_in(s[770]), .s(s[1033]), .c_out(c[1033]));
    fullAdder fa961 (.a(c[765]), .b(s[771]), .c_in(c[766]), .s(s[1034]), .c_out(c[1034]));
    fullAdder fa962 (.a(s[772]), .b(c[767]), .c_in(s[773]), .s(s[1035]), .c_out(c[1035]));
    fullAdder fa963 (.a(s[774]), .b(c[769]), .c_in(s[775]), .s(s[1036]), .c_out(c[1036]));
    fullAdder fa964 (.a(c[770]), .b(s[776]), .c_in(c[771]), .s(s[1037]), .c_out(c[1037]));
    fullAdder fa965 (.a(s[777]), .b(c[772]), .c_in(p[26][19]), .s(s[1038]), .c_out(c[1038]));
    fullAdder fa966 (.a(s[778]), .b(c[774]), .c_in(s[779]), .s(s[1039]), .c_out(c[1039]));
    fullAdder fa967 (.a(c[775]), .b(s[780]), .c_in(c[776]), .s(s[1040]), .c_out(c[1040]));
    halfAdder ha75 (.a(s[781]), .b(c[777]), .s(s[1041]), .c_out(c[1041]));
    fullAdder fa968 (.a(s[782]), .b(c[778]), .c_in(s[783]), .s(s[1042]), .c_out(c[1042]));
    fullAdder fa969 (.a(c[779]), .b(s[784]), .c_in(c[780]), .s(s[1043]), .c_out(c[1043]));
    halfAdder ha76 (.a(s[785]), .b(c[781]), .s(s[1044]), .c_out(c[1044]));
    fullAdder fa970 (.a(s[786]), .b(c[782]), .c_in(s[787]), .s(s[1045]), .c_out(c[1045]));
    fullAdder fa971 (.a(c[783]), .b(s[788]), .c_in(c[784]), .s(s[1046]), .c_out(c[1046]));
    halfAdder ha77 (.a(s[789]), .b(c[785]), .s(s[1047]), .c_out(c[1047]));
    fullAdder fa972 (.a(s[790]), .b(c[786]), .c_in(s[791]), .s(s[1048]), .c_out(c[1048]));
    fullAdder fa973 (.a(c[787]), .b(s[792]), .c_in(c[788]), .s(s[1049]), .c_out(c[1049]));
    halfAdder ha78 (.a(s[793]), .b(c[789]), .s(s[1050]), .c_out(c[1050]));
    fullAdder fa974 (.a(s[794]), .b(c[790]), .c_in(s[795]), .s(s[1051]), .c_out(c[1051]));
    fullAdder fa975 (.a(c[791]), .b(s[796]), .c_in(c[792]), .s(s[1052]), .c_out(c[1052]));
    halfAdder ha79 (.a(s[797]), .b(c[793]), .s(s[1053]), .c_out(c[1053]));
    fullAdder fa976 (.a(s[798]), .b(c[794]), .c_in(s[799]), .s(s[1054]), .c_out(c[1054]));
    fullAdder fa977 (.a(c[795]), .b(s[800]), .c_in(c[796]), .s(s[1055]), .c_out(c[1055]));
    halfAdder ha80 (.a(s[801]), .b(c[797]), .s(s[1056]), .c_out(c[1056]));
    fullAdder fa978 (.a(s[802]), .b(c[798]), .c_in(s[803]), .s(s[1057]), .c_out(c[1057]));
    fullAdder fa979 (.a(c[799]), .b(s[804]), .c_in(c[800]), .s(s[1058]), .c_out(c[1058]));
    halfAdder ha81 (.a(c[430]), .b(c[801]), .s(s[1059]), .c_out(c[1059]));
    fullAdder fa980 (.a(s[805]), .b(c[802]), .c_in(s[806]), .s(s[1060]), .c_out(c[1060]));
    fullAdder fa981 (.a(c[803]), .b(s[807]), .c_in(c[804]), .s(s[1061]), .c_out(c[1061]));
    fullAdder fa982 (.a(s[808]), .b(c[805]), .c_in(s[809]), .s(s[1062]), .c_out(c[1062]));
    fullAdder fa983 (.a(c[806]), .b(s[810]), .c_in(c[807]), .s(s[1063]), .c_out(c[1063]));
    fullAdder fa984 (.a(s[811]), .b(c[808]), .c_in(s[812]), .s(s[1064]), .c_out(c[1064]));
    fullAdder fa985 (.a(c[809]), .b(s[813]), .c_in(c[810]), .s(s[1065]), .c_out(c[1065]));
    fullAdder fa986 (.a(s[814]), .b(c[811]), .c_in(s[815]), .s(s[1066]), .c_out(c[1066]));
    fullAdder fa987 (.a(c[812]), .b(s[816]), .c_in(c[813]), .s(s[1067]), .c_out(c[1067]));
    fullAdder fa988 (.a(s[817]), .b(c[814]), .c_in(s[818]), .s(s[1068]), .c_out(c[1068]));
    fullAdder fa989 (.a(c[815]), .b(s[819]), .c_in(c[816]), .s(s[1069]), .c_out(c[1069]));
    fullAdder fa990 (.a(s[820]), .b(c[817]), .c_in(s[821]), .s(s[1070]), .c_out(c[1070]));
    fullAdder fa991 (.a(c[818]), .b(s[822]), .c_in(c[819]), .s(s[1071]), .c_out(c[1071]));
    fullAdder fa992 (.a(s[823]), .b(c[820]), .c_in(s[824]), .s(s[1072]), .c_out(c[1072]));
    fullAdder fa993 (.a(c[821]), .b(s[825]), .c_in(c[822]), .s(s[1073]), .c_out(c[1073]));
    fullAdder fa994 (.a(s[826]), .b(c[823]), .c_in(s[827]), .s(s[1074]), .c_out(c[1074]));
    fullAdder fa995 (.a(c[824]), .b(s[828]), .c_in(c[825]), .s(s[1075]), .c_out(c[1075]));
    fullAdder fa996 (.a(s[829]), .b(c[826]), .c_in(s[830]), .s(s[1076]), .c_out(c[1076]));
    fullAdder fa997 (.a(c[827]), .b(s[831]), .c_in(c[828]), .s(s[1077]), .c_out(c[1077]));
    fullAdder fa998 (.a(s[832]), .b(c[829]), .c_in(s[833]), .s(s[1078]), .c_out(c[1078]));
    fullAdder fa999 (.a(c[830]), .b(s[834]), .c_in(c[831]), .s(s[1079]), .c_out(c[1079]));
    fullAdder fa1000 (.a(s[835]), .b(c[832]), .c_in(s[836]), .s(s[1080]), .c_out(c[1080]));
    fullAdder fa1001 (.a(c[833]), .b(p[26][37]), .c_in(c[834]), .s(s[1081]), .c_out(c[1081]));
    fullAdder fa1002 (.a(s[837]), .b(c[835]), .c_in(s[838]), .s(s[1082]), .c_out(c[1082]));
    fullAdder fa1003 (.a(s[839]), .b(c[837]), .c_in(s[840]), .s(s[1083]), .c_out(c[1083]));
    fullAdder fa1004 (.a(s[841]), .b(c[839]), .c_in(s[842]), .s(s[1084]), .c_out(c[1084]));
    fullAdder fa1005 (.a(s[843]), .b(c[841]), .c_in(s[844]), .s(s[1085]), .c_out(c[1085]));
    fullAdder fa1006 (.a(s[845]), .b(c[843]), .c_in(s[846]), .s(s[1086]), .c_out(c[1086]));
    fullAdder fa1007 (.a(s[847]), .b(c[845]), .c_in(s[848]), .s(s[1087]), .c_out(c[1087]));
    fullAdder fa1008 (.a(s[849]), .b(c[847]), .c_in(c[496]), .s(s[1088]), .c_out(c[1088]));
    fullAdder fa1009 (.a(s[850]), .b(c[849]), .c_in(c[498]), .s(s[1089]), .c_out(c[1089]));
    fullAdder fa1010 (.a(s[851]), .b(c[850]), .c_in(c[500]), .s(s[1090]), .c_out(c[1090]));
    fullAdder fa1011 (.a(s[852]), .b(c[851]), .c_in(c[502]), .s(s[1091]), .c_out(c[1091]));
    fullAdder fa1012 (.a(s[853]), .b(c[852]), .c_in(c[504]), .s(s[1092]), .c_out(c[1092]));
    fullAdder fa1013 (.a(s[507]), .b(c[854]), .c_in(c[506]), .s(s[1093]), .c_out(c[1093]));
    fullAdder fa1014 (.a(1'b1), .b(c[855]), .c_in(p[26][53]), .s(s[1094]), .c_out(c[1094]));
    // Stage 4 Reduction
    fullAdder fa1015 (.a(s[2]), .b(c[856]), .c_in(c[1]), .s(s[1095]), .c_out(c[1095]));
    fullAdder fa1016 (.a(s[512]), .b(c[857]), .c_in(c[511]), .s(s[1096]), .c_out(c[1096]));
    fullAdder fa1017 (.a(s[860]), .b(c[859]), .c_in(c[515]), .s(s[1097]), .c_out(c[1097]));
    fullAdder fa1018 (.a(s[862]), .b(c[861]), .c_in(c[518]), .s(s[1098]), .c_out(c[1098]));
    fullAdder fa1019 (.a(s[863]), .b(c[862]), .c_in(c[520]), .s(s[1099]), .c_out(c[1099]));
    fullAdder fa1020 (.a(s[864]), .b(c[863]), .c_in(c[522]), .s(s[1100]), .c_out(c[1100]));
    fullAdder fa1021 (.a(s[865]), .b(c[864]), .c_in(s[866]), .s(s[1101]), .c_out(c[1101]));
    fullAdder fa1022 (.a(s[867]), .b(c[865]), .c_in(c[526]), .s(s[1102]), .c_out(c[1102]));
    fullAdder fa1023 (.a(s[868]), .b(c[867]), .c_in(s[869]), .s(s[1103]), .c_out(c[1103]));
    fullAdder fa1024 (.a(s[870]), .b(c[868]), .c_in(s[871]), .s(s[1104]), .c_out(c[1104]));
    fullAdder fa1025 (.a(s[872]), .b(c[870]), .c_in(s[873]), .s(s[1105]), .c_out(c[1105]));
    fullAdder fa1026 (.a(s[874]), .b(c[872]), .c_in(s[875]), .s(s[1106]), .c_out(c[1106]));
    fullAdder fa1027 (.a(s[876]), .b(c[874]), .c_in(s[877]), .s(s[1107]), .c_out(c[1107]));
    fullAdder fa1028 (.a(s[878]), .b(c[876]), .c_in(s[879]), .s(s[1108]), .c_out(c[1108]));
    fullAdder fa1029 (.a(s[880]), .b(c[878]), .c_in(s[881]), .s(s[1109]), .c_out(c[1109]));
    fullAdder fa1030 (.a(s[882]), .b(c[880]), .c_in(s[883]), .s(s[1110]), .c_out(c[1110]));
    fullAdder fa1031 (.a(s[884]), .b(c[882]), .c_in(s[885]), .s(s[1111]), .c_out(c[1111]));
    fullAdder fa1032 (.a(s[886]), .b(c[884]), .c_in(s[887]), .s(s[1112]), .c_out(c[1112]));
    fullAdder fa1033 (.a(s[888]), .b(c[886]), .c_in(s[889]), .s(s[1113]), .c_out(c[1113]));
    fullAdder fa1034 (.a(s[890]), .b(c[888]), .c_in(s[891]), .s(s[1114]), .c_out(c[1114]));
    fullAdder fa1035 (.a(s[893]), .b(c[890]), .c_in(s[894]), .s(s[1115]), .c_out(c[1115]));
    fullAdder fa1036 (.a(c[891]), .b(s[567]), .c_in(c[892]), .s(s[1116]), .c_out(c[1116]));
    fullAdder fa1037 (.a(s[895]), .b(c[893]), .c_in(s[896]), .s(s[1117]), .c_out(c[1117]));
    fullAdder fa1038 (.a(s[898]), .b(c[895]), .c_in(s[899]), .s(s[1118]), .c_out(c[1118]));
    fullAdder fa1039 (.a(c[896]), .b(s[900]), .c_in(c[897]), .s(s[1119]), .c_out(c[1119]));
    fullAdder fa1040 (.a(s[901]), .b(c[898]), .c_in(s[902]), .s(s[1120]), .c_out(c[1120]));
    fullAdder fa1041 (.a(c[899]), .b(s[903]), .c_in(c[900]), .s(s[1121]), .c_out(c[1121]));
    fullAdder fa1042 (.a(s[904]), .b(c[901]), .c_in(s[905]), .s(s[1122]), .c_out(c[1122]));
    fullAdder fa1043 (.a(c[902]), .b(s[906]), .c_in(c[903]), .s(s[1123]), .c_out(c[1123]));
    fullAdder fa1044 (.a(s[907]), .b(c[904]), .c_in(s[908]), .s(s[1124]), .c_out(c[1124]));
    fullAdder fa1045 (.a(c[905]), .b(s[909]), .c_in(c[906]), .s(s[1125]), .c_out(c[1125]));
    fullAdder fa1046 (.a(s[910]), .b(c[907]), .c_in(s[911]), .s(s[1126]), .c_out(c[1126]));
    fullAdder fa1047 (.a(c[908]), .b(s[912]), .c_in(c[909]), .s(s[1127]), .c_out(c[1127]));
    fullAdder fa1048 (.a(s[913]), .b(c[910]), .c_in(s[914]), .s(s[1128]), .c_out(c[1128]));
    fullAdder fa1049 (.a(c[911]), .b(s[915]), .c_in(c[912]), .s(s[1129]), .c_out(c[1129]));
    fullAdder fa1050 (.a(s[916]), .b(c[913]), .c_in(s[917]), .s(s[1130]), .c_out(c[1130]));
    fullAdder fa1051 (.a(c[914]), .b(s[918]), .c_in(c[915]), .s(s[1131]), .c_out(c[1131]));
    fullAdder fa1052 (.a(s[919]), .b(c[916]), .c_in(s[920]), .s(s[1132]), .c_out(c[1132]));
    fullAdder fa1053 (.a(c[917]), .b(s[921]), .c_in(c[918]), .s(s[1133]), .c_out(c[1133]));
    fullAdder fa1054 (.a(s[922]), .b(c[919]), .c_in(s[923]), .s(s[1134]), .c_out(c[1134]));
    fullAdder fa1055 (.a(c[920]), .b(s[924]), .c_in(c[921]), .s(s[1135]), .c_out(c[1135]));
    fullAdder fa1056 (.a(s[925]), .b(c[922]), .c_in(s[926]), .s(s[1136]), .c_out(c[1136]));
    fullAdder fa1057 (.a(c[923]), .b(s[927]), .c_in(c[924]), .s(s[1137]), .c_out(c[1137]));
    fullAdder fa1058 (.a(s[928]), .b(c[925]), .c_in(s[929]), .s(s[1138]), .c_out(c[1138]));
    fullAdder fa1059 (.a(c[926]), .b(s[930]), .c_in(c[927]), .s(s[1139]), .c_out(c[1139]));
    fullAdder fa1060 (.a(s[931]), .b(c[928]), .c_in(s[932]), .s(s[1140]), .c_out(c[1140]));
    fullAdder fa1061 (.a(c[929]), .b(s[933]), .c_in(c[930]), .s(s[1141]), .c_out(c[1141]));
    fullAdder fa1062 (.a(s[935]), .b(c[931]), .c_in(s[936]), .s(s[1142]), .c_out(c[1142]));
    fullAdder fa1063 (.a(c[932]), .b(s[937]), .c_in(c[933]), .s(s[1143]), .c_out(c[1143]));
    fullAdder fa1064 (.a(s[938]), .b(c[935]), .c_in(s[939]), .s(s[1144]), .c_out(c[1144]));
    fullAdder fa1065 (.a(c[936]), .b(s[940]), .c_in(c[937]), .s(s[1145]), .c_out(c[1145]));
    fullAdder fa1066 (.a(s[942]), .b(c[938]), .c_in(s[943]), .s(s[1146]), .c_out(c[1146]));
    fullAdder fa1067 (.a(c[939]), .b(s[944]), .c_in(c[940]), .s(s[1147]), .c_out(c[1147]));
    fullAdder fa1068 (.a(s[946]), .b(c[942]), .c_in(s[947]), .s(s[1148]), .c_out(c[1148]));
    fullAdder fa1069 (.a(c[943]), .b(s[948]), .c_in(c[944]), .s(s[1149]), .c_out(c[1149]));
    fullAdder fa1070 (.a(s[950]), .b(c[946]), .c_in(s[951]), .s(s[1150]), .c_out(c[1150]));
    fullAdder fa1071 (.a(c[947]), .b(s[952]), .c_in(c[948]), .s(s[1151]), .c_out(c[1151]));
    fullAdder fa1072 (.a(s[954]), .b(c[950]), .c_in(s[955]), .s(s[1152]), .c_out(c[1152]));
    fullAdder fa1073 (.a(c[951]), .b(s[956]), .c_in(c[952]), .s(s[1153]), .c_out(c[1153]));
    fullAdder fa1074 (.a(s[958]), .b(c[954]), .c_in(s[959]), .s(s[1154]), .c_out(c[1154]));
    fullAdder fa1075 (.a(c[955]), .b(s[960]), .c_in(c[956]), .s(s[1155]), .c_out(c[1155]));
    fullAdder fa1076 (.a(s[962]), .b(c[958]), .c_in(s[963]), .s(s[1156]), .c_out(c[1156]));
    fullAdder fa1077 (.a(c[959]), .b(s[964]), .c_in(c[960]), .s(s[1157]), .c_out(c[1157]));
    fullAdder fa1078 (.a(s[966]), .b(c[962]), .c_in(s[967]), .s(s[1158]), .c_out(c[1158]));
    fullAdder fa1079 (.a(c[963]), .b(s[968]), .c_in(c[964]), .s(s[1159]), .c_out(c[1159]));
    fullAdder fa1080 (.a(s[970]), .b(c[966]), .c_in(s[971]), .s(s[1160]), .c_out(c[1160]));
    fullAdder fa1081 (.a(c[967]), .b(s[972]), .c_in(c[968]), .s(s[1161]), .c_out(c[1161]));
    fullAdder fa1082 (.a(s[974]), .b(c[970]), .c_in(s[975]), .s(s[1162]), .c_out(c[1162]));
    fullAdder fa1083 (.a(c[971]), .b(s[976]), .c_in(c[972]), .s(s[1163]), .c_out(c[1163]));
    fullAdder fa1084 (.a(s[978]), .b(c[974]), .c_in(s[979]), .s(s[1164]), .c_out(c[1164]));
    fullAdder fa1085 (.a(c[975]), .b(s[980]), .c_in(c[976]), .s(s[1165]), .c_out(c[1165]));
    fullAdder fa1086 (.a(s[982]), .b(c[978]), .c_in(s[983]), .s(s[1166]), .c_out(c[1166]));
    fullAdder fa1087 (.a(c[979]), .b(s[984]), .c_in(c[980]), .s(s[1167]), .c_out(c[1167]));
    fullAdder fa1088 (.a(s[986]), .b(c[982]), .c_in(s[987]), .s(s[1168]), .c_out(c[1168]));
    fullAdder fa1089 (.a(c[983]), .b(s[988]), .c_in(c[984]), .s(s[1169]), .c_out(c[1169]));
    fullAdder fa1090 (.a(s[990]), .b(c[986]), .c_in(s[991]), .s(s[1170]), .c_out(c[1170]));
    fullAdder fa1091 (.a(c[987]), .b(s[992]), .c_in(c[988]), .s(s[1171]), .c_out(c[1171]));
    fullAdder fa1092 (.a(s[994]), .b(c[990]), .c_in(s[995]), .s(s[1172]), .c_out(c[1172]));
    fullAdder fa1093 (.a(c[991]), .b(s[996]), .c_in(c[992]), .s(s[1173]), .c_out(c[1173]));
    fullAdder fa1094 (.a(s[998]), .b(c[994]), .c_in(s[999]), .s(s[1174]), .c_out(c[1174]));
    fullAdder fa1095 (.a(c[995]), .b(s[1000]), .c_in(c[996]), .s(s[1175]), .c_out(c[1175]));
    fullAdder fa1096 (.a(s[1002]), .b(c[998]), .c_in(s[1003]), .s(s[1176]), .c_out(c[1176]));
    fullAdder fa1097 (.a(c[999]), .b(s[1004]), .c_in(c[1000]), .s(s[1177]), .c_out(c[1177]));
    fullAdder fa1098 (.a(s[1006]), .b(c[1002]), .c_in(s[1007]), .s(s[1178]), .c_out(c[1178]));
    fullAdder fa1099 (.a(c[1003]), .b(s[1008]), .c_in(c[1004]), .s(s[1179]), .c_out(c[1179]));
    fullAdder fa1100 (.a(s[1010]), .b(c[1006]), .c_in(s[1011]), .s(s[1180]), .c_out(c[1180]));
    fullAdder fa1101 (.a(c[1007]), .b(s[1012]), .c_in(c[1008]), .s(s[1181]), .c_out(c[1181]));
    fullAdder fa1102 (.a(s[1014]), .b(c[1010]), .c_in(s[1015]), .s(s[1182]), .c_out(c[1182]));
    fullAdder fa1103 (.a(c[1011]), .b(s[1016]), .c_in(c[1012]), .s(s[1183]), .c_out(c[1183]));
    fullAdder fa1104 (.a(s[1018]), .b(c[1014]), .c_in(s[1019]), .s(s[1184]), .c_out(c[1184]));
    fullAdder fa1105 (.a(c[1015]), .b(s[1020]), .c_in(c[1016]), .s(s[1185]), .c_out(c[1185]));
    fullAdder fa1106 (.a(s[1021]), .b(c[1018]), .c_in(s[1022]), .s(s[1186]), .c_out(c[1186]));
    fullAdder fa1107 (.a(c[1019]), .b(s[1023]), .c_in(c[1020]), .s(s[1187]), .c_out(c[1187]));
    fullAdder fa1108 (.a(s[1024]), .b(c[1021]), .c_in(s[1025]), .s(s[1188]), .c_out(c[1188]));
    fullAdder fa1109 (.a(c[1022]), .b(s[1026]), .c_in(c[1023]), .s(s[1189]), .c_out(c[1189]));
    fullAdder fa1110 (.a(s[1027]), .b(c[1024]), .c_in(s[1028]), .s(s[1190]), .c_out(c[1190]));
    fullAdder fa1111 (.a(c[1025]), .b(s[1029]), .c_in(c[1026]), .s(s[1191]), .c_out(c[1191]));
    fullAdder fa1112 (.a(s[1030]), .b(c[1027]), .c_in(s[1031]), .s(s[1192]), .c_out(c[1192]));
    fullAdder fa1113 (.a(c[1028]), .b(s[1032]), .c_in(c[1029]), .s(s[1193]), .c_out(c[1193]));
    fullAdder fa1114 (.a(s[1033]), .b(c[1030]), .c_in(s[1034]), .s(s[1194]), .c_out(c[1194]));
    fullAdder fa1115 (.a(c[1031]), .b(s[1035]), .c_in(c[1032]), .s(s[1195]), .c_out(c[1195]));
    fullAdder fa1116 (.a(s[1036]), .b(c[1033]), .c_in(s[1037]), .s(s[1196]), .c_out(c[1196]));
    fullAdder fa1117 (.a(c[1034]), .b(s[1038]), .c_in(c[1035]), .s(s[1197]), .c_out(c[1197]));
    fullAdder fa1118 (.a(s[1039]), .b(c[1036]), .c_in(s[1040]), .s(s[1198]), .c_out(c[1198]));
    fullAdder fa1119 (.a(c[1037]), .b(s[1041]), .c_in(c[1038]), .s(s[1199]), .c_out(c[1199]));
    fullAdder fa1120 (.a(s[1042]), .b(c[1039]), .c_in(s[1043]), .s(s[1200]), .c_out(c[1200]));
    fullAdder fa1121 (.a(c[1040]), .b(s[1044]), .c_in(c[1041]), .s(s[1201]), .c_out(c[1201]));
    fullAdder fa1122 (.a(s[1045]), .b(c[1042]), .c_in(s[1046]), .s(s[1202]), .c_out(c[1202]));
    fullAdder fa1123 (.a(c[1043]), .b(s[1047]), .c_in(c[1044]), .s(s[1203]), .c_out(c[1203]));
    fullAdder fa1124 (.a(s[1048]), .b(c[1045]), .c_in(s[1049]), .s(s[1204]), .c_out(c[1204]));
    fullAdder fa1125 (.a(c[1046]), .b(s[1050]), .c_in(c[1047]), .s(s[1205]), .c_out(c[1205]));
    fullAdder fa1126 (.a(s[1051]), .b(c[1048]), .c_in(s[1052]), .s(s[1206]), .c_out(c[1206]));
    fullAdder fa1127 (.a(c[1049]), .b(s[1053]), .c_in(c[1050]), .s(s[1207]), .c_out(c[1207]));
    fullAdder fa1128 (.a(s[1054]), .b(c[1051]), .c_in(s[1055]), .s(s[1208]), .c_out(c[1208]));
    fullAdder fa1129 (.a(c[1052]), .b(s[1056]), .c_in(c[1053]), .s(s[1209]), .c_out(c[1209]));
    fullAdder fa1130 (.a(s[1057]), .b(c[1054]), .c_in(s[1058]), .s(s[1210]), .c_out(c[1210]));
    fullAdder fa1131 (.a(c[1055]), .b(s[1059]), .c_in(c[1056]), .s(s[1211]), .c_out(c[1211]));
    fullAdder fa1132 (.a(s[1060]), .b(c[1057]), .c_in(s[1061]), .s(s[1212]), .c_out(c[1212]));
    fullAdder fa1133 (.a(c[1058]), .b(c[435]), .c_in(c[1059]), .s(s[1213]), .c_out(c[1213]));
    fullAdder fa1134 (.a(s[1062]), .b(c[1060]), .c_in(s[1063]), .s(s[1214]), .c_out(c[1214]));
    fullAdder fa1135 (.a(s[1064]), .b(c[1062]), .c_in(s[1065]), .s(s[1215]), .c_out(c[1215]));
    fullAdder fa1136 (.a(s[1066]), .b(c[1064]), .c_in(s[1067]), .s(s[1216]), .c_out(c[1216]));
    fullAdder fa1137 (.a(s[1068]), .b(c[1066]), .c_in(s[1069]), .s(s[1217]), .c_out(c[1217]));
    fullAdder fa1138 (.a(s[1070]), .b(c[1068]), .c_in(s[1071]), .s(s[1218]), .c_out(c[1218]));
    fullAdder fa1139 (.a(s[1072]), .b(c[1070]), .c_in(s[1073]), .s(s[1219]), .c_out(c[1219]));
    fullAdder fa1140 (.a(s[1074]), .b(c[1072]), .c_in(s[1075]), .s(s[1220]), .c_out(c[1220]));
    fullAdder fa1141 (.a(s[1076]), .b(c[1074]), .c_in(s[1077]), .s(s[1221]), .c_out(c[1221]));
    fullAdder fa1142 (.a(s[1078]), .b(c[1076]), .c_in(s[1079]), .s(s[1222]), .c_out(c[1222]));
    fullAdder fa1143 (.a(s[1080]), .b(c[1078]), .c_in(s[1081]), .s(s[1223]), .c_out(c[1223]));
    fullAdder fa1144 (.a(s[1082]), .b(c[1080]), .c_in(c[836]), .s(s[1224]), .c_out(c[1224]));
    fullAdder fa1145 (.a(s[1083]), .b(c[1082]), .c_in(c[838]), .s(s[1225]), .c_out(c[1225]));
    fullAdder fa1146 (.a(s[1084]), .b(c[1083]), .c_in(c[840]), .s(s[1226]), .c_out(c[1226]));
    fullAdder fa1147 (.a(s[1085]), .b(c[1084]), .c_in(c[842]), .s(s[1227]), .c_out(c[1227]));
    fullAdder fa1148 (.a(s[1086]), .b(c[1085]), .c_in(c[844]), .s(s[1228]), .c_out(c[1228]));
    fullAdder fa1149 (.a(s[1087]), .b(c[1086]), .c_in(c[846]), .s(s[1229]), .c_out(c[1229]));
    fullAdder fa1150 (.a(s[1088]), .b(c[1087]), .c_in(c[848]), .s(s[1230]), .c_out(c[1230]));
    fullAdder fa1151 (.a(s[854]), .b(c[1092]), .c_in(c[853]), .s(s[1231]), .c_out(c[1231]));
    fullAdder fa1152 (.a(s[508]), .b(c[1093]), .c_in(c[507]), .s(s[1232]), .c_out(c[1232]));
    // Stage 5 Reduction
    fullAdder fa1153 (.a(s[861]), .b(c[1097]), .c_in(c[860]), .s(s[1233]), .c_out(c[1233]));
    fullAdder fa1154 (.a(s[1102]), .b(c[1101]), .c_in(c[866]), .s(s[1234]), .c_out(c[1234]));
    fullAdder fa1155 (.a(s[1104]), .b(c[1103]), .c_in(c[869]), .s(s[1235]), .c_out(c[1235]));
    fullAdder fa1156 (.a(s[1105]), .b(c[1104]), .c_in(c[871]), .s(s[1236]), .c_out(c[1236]));
    fullAdder fa1157 (.a(s[1106]), .b(c[1105]), .c_in(c[873]), .s(s[1237]), .c_out(c[1237]));
    fullAdder fa1158 (.a(s[1107]), .b(c[1106]), .c_in(c[875]), .s(s[1238]), .c_out(c[1238]));
    fullAdder fa1159 (.a(s[1108]), .b(c[1107]), .c_in(c[877]), .s(s[1239]), .c_out(c[1239]));
    fullAdder fa1160 (.a(s[1109]), .b(c[1108]), .c_in(c[879]), .s(s[1240]), .c_out(c[1240]));
    fullAdder fa1161 (.a(s[1110]), .b(c[1109]), .c_in(c[881]), .s(s[1241]), .c_out(c[1241]));
    fullAdder fa1162 (.a(s[1111]), .b(c[1110]), .c_in(c[883]), .s(s[1242]), .c_out(c[1242]));
    fullAdder fa1163 (.a(s[1112]), .b(c[1111]), .c_in(c[885]), .s(s[1243]), .c_out(c[1243]));
    fullAdder fa1164 (.a(s[1113]), .b(c[1112]), .c_in(c[887]), .s(s[1244]), .c_out(c[1244]));
    fullAdder fa1165 (.a(s[1114]), .b(c[1113]), .c_in(c[889]), .s(s[1245]), .c_out(c[1245]));
    fullAdder fa1166 (.a(s[1115]), .b(c[1114]), .c_in(s[1116]), .s(s[1246]), .c_out(c[1246]));
    fullAdder fa1167 (.a(s[1117]), .b(c[1115]), .c_in(c[894]), .s(s[1247]), .c_out(c[1247]));
    halfAdder ha82 (.a(c[1116]), .b(s[897]), .s(s[1248]), .c_out(c[1248]));
    fullAdder fa1168 (.a(s[1118]), .b(c[1117]), .c_in(s[1119]), .s(s[1249]), .c_out(c[1249]));
    fullAdder fa1169 (.a(s[1120]), .b(c[1118]), .c_in(s[1121]), .s(s[1250]), .c_out(c[1250]));
    fullAdder fa1170 (.a(s[1122]), .b(c[1120]), .c_in(s[1123]), .s(s[1251]), .c_out(c[1251]));
    fullAdder fa1171 (.a(s[1124]), .b(c[1122]), .c_in(s[1125]), .s(s[1252]), .c_out(c[1252]));
    fullAdder fa1172 (.a(s[1126]), .b(c[1124]), .c_in(s[1127]), .s(s[1253]), .c_out(c[1253]));
    fullAdder fa1173 (.a(s[1128]), .b(c[1126]), .c_in(s[1129]), .s(s[1254]), .c_out(c[1254]));
    fullAdder fa1174 (.a(s[1130]), .b(c[1128]), .c_in(s[1131]), .s(s[1255]), .c_out(c[1255]));
    halfAdder ha83 (.a(c[1129]), .b(c[596]), .s(s[1256]), .c_out(c[1256]));
    fullAdder fa1175 (.a(s[1132]), .b(c[1130]), .c_in(s[1133]), .s(s[1257]), .c_out(c[1257]));
    fullAdder fa1176 (.a(s[1134]), .b(c[1132]), .c_in(s[1135]), .s(s[1258]), .c_out(c[1258]));
    halfAdder ha84 (.a(c[1133]), .b(c[605]), .s(s[1259]), .c_out(c[1259]));
    fullAdder fa1177 (.a(s[1136]), .b(c[1134]), .c_in(s[1137]), .s(s[1260]), .c_out(c[1260]));
    halfAdder ha85 (.a(c[1135]), .b(c[610]), .s(s[1261]), .c_out(c[1261]));
    fullAdder fa1178 (.a(s[1138]), .b(c[1136]), .c_in(s[1139]), .s(s[1262]), .c_out(c[1262]));
    halfAdder ha86 (.a(c[1137]), .b(c[615]), .s(s[1263]), .c_out(c[1263]));
    fullAdder fa1179 (.a(s[1140]), .b(c[1138]), .c_in(s[1141]), .s(s[1264]), .c_out(c[1264]));
    halfAdder ha87 (.a(c[1139]), .b(s[934]), .s(s[1265]), .c_out(c[1265]));
    fullAdder fa1180 (.a(s[1142]), .b(c[1140]), .c_in(s[1143]), .s(s[1266]), .c_out(c[1266]));
    fullAdder fa1181 (.a(c[1141]), .b(c[625]), .c_in(c[934]), .s(s[1267]), .c_out(c[1267]));
    fullAdder fa1182 (.a(s[1144]), .b(c[1142]), .c_in(s[1145]), .s(s[1268]), .c_out(c[1268]));
    halfAdder ha88 (.a(c[1143]), .b(s[941]), .s(s[1269]), .c_out(c[1269]));
    fullAdder fa1183 (.a(s[1146]), .b(c[1144]), .c_in(s[1147]), .s(s[1270]), .c_out(c[1270]));
    fullAdder fa1184 (.a(c[1145]), .b(s[945]), .c_in(c[941]), .s(s[1271]), .c_out(c[1271]));
    fullAdder fa1185 (.a(s[1148]), .b(c[1146]), .c_in(s[1149]), .s(s[1272]), .c_out(c[1272]));
    fullAdder fa1186 (.a(c[1147]), .b(s[949]), .c_in(c[945]), .s(s[1273]), .c_out(c[1273]));
    fullAdder fa1187 (.a(s[1150]), .b(c[1148]), .c_in(s[1151]), .s(s[1274]), .c_out(c[1274]));
    fullAdder fa1188 (.a(c[1149]), .b(s[953]), .c_in(c[949]), .s(s[1275]), .c_out(c[1275]));
    fullAdder fa1189 (.a(s[1152]), .b(c[1150]), .c_in(s[1153]), .s(s[1276]), .c_out(c[1276]));
    fullAdder fa1190 (.a(c[1151]), .b(s[957]), .c_in(c[953]), .s(s[1277]), .c_out(c[1277]));
    fullAdder fa1191 (.a(s[1154]), .b(c[1152]), .c_in(s[1155]), .s(s[1278]), .c_out(c[1278]));
    fullAdder fa1192 (.a(c[1153]), .b(s[961]), .c_in(c[957]), .s(s[1279]), .c_out(c[1279]));
    fullAdder fa1193 (.a(s[1156]), .b(c[1154]), .c_in(s[1157]), .s(s[1280]), .c_out(c[1280]));
    fullAdder fa1194 (.a(c[1155]), .b(s[965]), .c_in(c[961]), .s(s[1281]), .c_out(c[1281]));
    fullAdder fa1195 (.a(s[1158]), .b(c[1156]), .c_in(s[1159]), .s(s[1282]), .c_out(c[1282]));
    fullAdder fa1196 (.a(c[1157]), .b(s[969]), .c_in(c[965]), .s(s[1283]), .c_out(c[1283]));
    fullAdder fa1197 (.a(s[1160]), .b(c[1158]), .c_in(s[1161]), .s(s[1284]), .c_out(c[1284]));
    fullAdder fa1198 (.a(c[1159]), .b(s[973]), .c_in(c[969]), .s(s[1285]), .c_out(c[1285]));
    fullAdder fa1199 (.a(s[1162]), .b(c[1160]), .c_in(s[1163]), .s(s[1286]), .c_out(c[1286]));
    fullAdder fa1200 (.a(c[1161]), .b(s[977]), .c_in(c[973]), .s(s[1287]), .c_out(c[1287]));
    fullAdder fa1201 (.a(s[1164]), .b(c[1162]), .c_in(s[1165]), .s(s[1288]), .c_out(c[1288]));
    fullAdder fa1202 (.a(c[1163]), .b(s[981]), .c_in(c[977]), .s(s[1289]), .c_out(c[1289]));
    fullAdder fa1203 (.a(s[1166]), .b(c[1164]), .c_in(s[1167]), .s(s[1290]), .c_out(c[1290]));
    fullAdder fa1204 (.a(c[1165]), .b(s[985]), .c_in(c[981]), .s(s[1291]), .c_out(c[1291]));
    fullAdder fa1205 (.a(s[1168]), .b(c[1166]), .c_in(s[1169]), .s(s[1292]), .c_out(c[1292]));
    fullAdder fa1206 (.a(c[1167]), .b(s[989]), .c_in(c[985]), .s(s[1293]), .c_out(c[1293]));
    fullAdder fa1207 (.a(s[1170]), .b(c[1168]), .c_in(s[1171]), .s(s[1294]), .c_out(c[1294]));
    fullAdder fa1208 (.a(c[1169]), .b(s[993]), .c_in(c[989]), .s(s[1295]), .c_out(c[1295]));
    fullAdder fa1209 (.a(s[1172]), .b(c[1170]), .c_in(s[1173]), .s(s[1296]), .c_out(c[1296]));
    fullAdder fa1210 (.a(c[1171]), .b(s[997]), .c_in(c[993]), .s(s[1297]), .c_out(c[1297]));
    fullAdder fa1211 (.a(s[1174]), .b(c[1172]), .c_in(s[1175]), .s(s[1298]), .c_out(c[1298]));
    fullAdder fa1212 (.a(c[1173]), .b(s[1001]), .c_in(c[997]), .s(s[1299]), .c_out(c[1299]));
    fullAdder fa1213 (.a(s[1176]), .b(c[1174]), .c_in(s[1177]), .s(s[1300]), .c_out(c[1300]));
    fullAdder fa1214 (.a(c[1175]), .b(s[1005]), .c_in(c[1001]), .s(s[1301]), .c_out(c[1301]));
    fullAdder fa1215 (.a(s[1178]), .b(c[1176]), .c_in(s[1179]), .s(s[1302]), .c_out(c[1302]));
    fullAdder fa1216 (.a(c[1177]), .b(s[1009]), .c_in(c[1005]), .s(s[1303]), .c_out(c[1303]));
    fullAdder fa1217 (.a(s[1180]), .b(c[1178]), .c_in(s[1181]), .s(s[1304]), .c_out(c[1304]));
    fullAdder fa1218 (.a(c[1179]), .b(s[1013]), .c_in(c[1009]), .s(s[1305]), .c_out(c[1305]));
    fullAdder fa1219 (.a(s[1182]), .b(c[1180]), .c_in(s[1183]), .s(s[1306]), .c_out(c[1306]));
    fullAdder fa1220 (.a(c[1181]), .b(s[1017]), .c_in(c[1013]), .s(s[1307]), .c_out(c[1307]));
    fullAdder fa1221 (.a(s[1184]), .b(c[1182]), .c_in(s[1185]), .s(s[1308]), .c_out(c[1308]));
    fullAdder fa1222 (.a(c[1183]), .b(c[743]), .c_in(c[1017]), .s(s[1309]), .c_out(c[1309]));
    fullAdder fa1223 (.a(s[1186]), .b(c[1184]), .c_in(s[1187]), .s(s[1310]), .c_out(c[1310]));
    halfAdder ha89 (.a(c[1185]), .b(c[748]), .s(s[1311]), .c_out(c[1311]));
    fullAdder fa1224 (.a(s[1188]), .b(c[1186]), .c_in(s[1189]), .s(s[1312]), .c_out(c[1312]));
    halfAdder ha90 (.a(c[1187]), .b(c[753]), .s(s[1313]), .c_out(c[1313]));
    fullAdder fa1225 (.a(s[1190]), .b(c[1188]), .c_in(s[1191]), .s(s[1314]), .c_out(c[1314]));
    halfAdder ha91 (.a(c[1189]), .b(c[758]), .s(s[1315]), .c_out(c[1315]));
    fullAdder fa1226 (.a(s[1192]), .b(c[1190]), .c_in(s[1193]), .s(s[1316]), .c_out(c[1316]));
    halfAdder ha92 (.a(c[1191]), .b(c[763]), .s(s[1317]), .c_out(c[1317]));
    fullAdder fa1227 (.a(s[1194]), .b(c[1192]), .c_in(s[1195]), .s(s[1318]), .c_out(c[1318]));
    halfAdder ha93 (.a(c[1193]), .b(c[768]), .s(s[1319]), .c_out(c[1319]));
    fullAdder fa1228 (.a(s[1196]), .b(c[1194]), .c_in(s[1197]), .s(s[1320]), .c_out(c[1320]));
    halfAdder ha94 (.a(c[1195]), .b(c[773]), .s(s[1321]), .c_out(c[1321]));
    fullAdder fa1229 (.a(s[1198]), .b(c[1196]), .c_in(s[1199]), .s(s[1322]), .c_out(c[1322]));
    fullAdder fa1230 (.a(s[1200]), .b(c[1198]), .c_in(s[1201]), .s(s[1323]), .c_out(c[1323]));
    fullAdder fa1231 (.a(s[1202]), .b(c[1200]), .c_in(s[1203]), .s(s[1324]), .c_out(c[1324]));
    fullAdder fa1232 (.a(s[1204]), .b(c[1202]), .c_in(s[1205]), .s(s[1325]), .c_out(c[1325]));
    fullAdder fa1233 (.a(s[1206]), .b(c[1204]), .c_in(s[1207]), .s(s[1326]), .c_out(c[1326]));
    fullAdder fa1234 (.a(s[1208]), .b(c[1206]), .c_in(s[1209]), .s(s[1327]), .c_out(c[1327]));
    fullAdder fa1235 (.a(s[1210]), .b(c[1208]), .c_in(s[1211]), .s(s[1328]), .c_out(c[1328]));
    fullAdder fa1236 (.a(s[1212]), .b(c[1210]), .c_in(s[1213]), .s(s[1329]), .c_out(c[1329]));
    fullAdder fa1237 (.a(s[1214]), .b(c[1212]), .c_in(c[1061]), .s(s[1330]), .c_out(c[1330]));
    halfAdder ha95 (.a(c[1213]), .b(c[440]), .s(s[1331]), .c_out(c[1331]));
    fullAdder fa1238 (.a(s[1215]), .b(c[1214]), .c_in(c[1063]), .s(s[1332]), .c_out(c[1332]));
    fullAdder fa1239 (.a(s[1216]), .b(c[1215]), .c_in(c[1065]), .s(s[1333]), .c_out(c[1333]));
    fullAdder fa1240 (.a(s[1217]), .b(c[1216]), .c_in(c[1067]), .s(s[1334]), .c_out(c[1334]));
    fullAdder fa1241 (.a(s[1218]), .b(c[1217]), .c_in(c[1069]), .s(s[1335]), .c_out(c[1335]));
    fullAdder fa1242 (.a(s[1219]), .b(c[1218]), .c_in(c[1071]), .s(s[1336]), .c_out(c[1336]));
    fullAdder fa1243 (.a(s[1220]), .b(c[1219]), .c_in(c[1073]), .s(s[1337]), .c_out(c[1337]));
    fullAdder fa1244 (.a(s[1221]), .b(c[1220]), .c_in(c[1075]), .s(s[1338]), .c_out(c[1338]));
    fullAdder fa1245 (.a(s[1222]), .b(c[1221]), .c_in(c[1077]), .s(s[1339]), .c_out(c[1339]));
    fullAdder fa1246 (.a(s[1223]), .b(c[1222]), .c_in(c[1079]), .s(s[1340]), .c_out(c[1340]));
    fullAdder fa1247 (.a(s[1224]), .b(c[1223]), .c_in(c[1081]), .s(s[1341]), .c_out(c[1341]));
    fullAdder fa1248 (.a(s[1089]), .b(c[1230]), .c_in(c[1088]), .s(s[1342]), .c_out(c[1342]));
    // Stage 6 Reduction
    fullAdder fa1249 (.a(s[1103]), .b(c[1234]), .c_in(c[1102]), .s(s[1343]), .c_out(c[1343]));
    fullAdder fa1250 (.a(s[1241]), .b(c[1240]), .c_in(c[58]), .s(s[1344]), .c_out(c[1344]));
    fullAdder fa1251 (.a(s[1243]), .b(c[1242]), .c_in(c[67]), .s(s[1345]), .c_out(c[1345]));
    fullAdder fa1252 (.a(s[1244]), .b(c[1243]), .c_in(s[560]), .s(s[1346]), .c_out(c[1346]));
    fullAdder fa1253 (.a(s[1245]), .b(c[1244]), .c_in(s[892]), .s(s[1347]), .c_out(c[1347]));
    fullAdder fa1254 (.a(s[1247]), .b(c[1246]), .c_in(s[1248]), .s(s[1348]), .c_out(c[1348]));
    fullAdder fa1255 (.a(s[1249]), .b(c[1247]), .c_in(c[1248]), .s(s[1349]), .c_out(c[1349]));
    fullAdder fa1256 (.a(s[1250]), .b(c[1249]), .c_in(c[1119]), .s(s[1350]), .c_out(c[1350]));
    fullAdder fa1257 (.a(s[1251]), .b(c[1250]), .c_in(c[1121]), .s(s[1351]), .c_out(c[1351]));
    fullAdder fa1258 (.a(s[1252]), .b(c[1251]), .c_in(c[1123]), .s(s[1352]), .c_out(c[1352]));
    fullAdder fa1259 (.a(s[1253]), .b(c[1252]), .c_in(c[1125]), .s(s[1353]), .c_out(c[1353]));
    fullAdder fa1260 (.a(s[1254]), .b(c[1253]), .c_in(c[1127]), .s(s[1354]), .c_out(c[1354]));
    fullAdder fa1261 (.a(s[1255]), .b(c[1254]), .c_in(s[1256]), .s(s[1355]), .c_out(c[1355]));
    fullAdder fa1262 (.a(s[1257]), .b(c[1255]), .c_in(c[1131]), .s(s[1356]), .c_out(c[1356]));
    fullAdder fa1263 (.a(s[1258]), .b(c[1257]), .c_in(s[1259]), .s(s[1357]), .c_out(c[1357]));
    fullAdder fa1264 (.a(s[1260]), .b(c[1258]), .c_in(s[1261]), .s(s[1358]), .c_out(c[1358]));
    fullAdder fa1265 (.a(s[1262]), .b(c[1260]), .c_in(s[1263]), .s(s[1359]), .c_out(c[1359]));
    fullAdder fa1266 (.a(s[1264]), .b(c[1262]), .c_in(s[1265]), .s(s[1360]), .c_out(c[1360]));
    fullAdder fa1267 (.a(s[1266]), .b(c[1264]), .c_in(s[1267]), .s(s[1361]), .c_out(c[1361]));
    fullAdder fa1268 (.a(s[1268]), .b(c[1266]), .c_in(s[1269]), .s(s[1362]), .c_out(c[1362]));
    fullAdder fa1269 (.a(s[1270]), .b(c[1268]), .c_in(s[1271]), .s(s[1363]), .c_out(c[1363]));
    fullAdder fa1270 (.a(s[1272]), .b(c[1270]), .c_in(s[1273]), .s(s[1364]), .c_out(c[1364]));
    fullAdder fa1271 (.a(s[1274]), .b(c[1272]), .c_in(s[1275]), .s(s[1365]), .c_out(c[1365]));
    fullAdder fa1272 (.a(s[1276]), .b(c[1274]), .c_in(s[1277]), .s(s[1366]), .c_out(c[1366]));
    fullAdder fa1273 (.a(s[1278]), .b(c[1276]), .c_in(s[1279]), .s(s[1367]), .c_out(c[1367]));
    fullAdder fa1274 (.a(s[1280]), .b(c[1278]), .c_in(s[1281]), .s(s[1368]), .c_out(c[1368]));
    fullAdder fa1275 (.a(s[1282]), .b(c[1280]), .c_in(s[1283]), .s(s[1369]), .c_out(c[1369]));
    fullAdder fa1276 (.a(s[1284]), .b(c[1282]), .c_in(s[1285]), .s(s[1370]), .c_out(c[1370]));
    fullAdder fa1277 (.a(s[1286]), .b(c[1284]), .c_in(s[1287]), .s(s[1371]), .c_out(c[1371]));
    fullAdder fa1278 (.a(s[1288]), .b(c[1286]), .c_in(s[1289]), .s(s[1372]), .c_out(c[1372]));
    fullAdder fa1279 (.a(s[1290]), .b(c[1288]), .c_in(s[1291]), .s(s[1373]), .c_out(c[1373]));
    fullAdder fa1280 (.a(s[1292]), .b(c[1290]), .c_in(s[1293]), .s(s[1374]), .c_out(c[1374]));
    fullAdder fa1281 (.a(s[1294]), .b(c[1292]), .c_in(s[1295]), .s(s[1375]), .c_out(c[1375]));
    fullAdder fa1282 (.a(s[1296]), .b(c[1294]), .c_in(s[1297]), .s(s[1376]), .c_out(c[1376]));
    fullAdder fa1283 (.a(s[1298]), .b(c[1296]), .c_in(s[1299]), .s(s[1377]), .c_out(c[1377]));
    fullAdder fa1284 (.a(s[1300]), .b(c[1298]), .c_in(s[1301]), .s(s[1378]), .c_out(c[1378]));
    fullAdder fa1285 (.a(s[1302]), .b(c[1300]), .c_in(s[1303]), .s(s[1379]), .c_out(c[1379]));
    fullAdder fa1286 (.a(s[1304]), .b(c[1302]), .c_in(s[1305]), .s(s[1380]), .c_out(c[1380]));
    fullAdder fa1287 (.a(s[1306]), .b(c[1304]), .c_in(s[1307]), .s(s[1381]), .c_out(c[1381]));
    fullAdder fa1288 (.a(s[1308]), .b(c[1306]), .c_in(s[1309]), .s(s[1382]), .c_out(c[1382]));
    fullAdder fa1289 (.a(s[1310]), .b(c[1308]), .c_in(s[1311]), .s(s[1383]), .c_out(c[1383]));
    fullAdder fa1290 (.a(s[1312]), .b(c[1310]), .c_in(s[1313]), .s(s[1384]), .c_out(c[1384]));
    fullAdder fa1291 (.a(s[1314]), .b(c[1312]), .c_in(s[1315]), .s(s[1385]), .c_out(c[1385]));
    fullAdder fa1292 (.a(s[1316]), .b(c[1314]), .c_in(s[1317]), .s(s[1386]), .c_out(c[1386]));
    fullAdder fa1293 (.a(s[1318]), .b(c[1316]), .c_in(s[1319]), .s(s[1387]), .c_out(c[1387]));
    fullAdder fa1294 (.a(s[1320]), .b(c[1318]), .c_in(s[1321]), .s(s[1388]), .c_out(c[1388]));
    fullAdder fa1295 (.a(s[1322]), .b(c[1320]), .c_in(c[1197]), .s(s[1389]), .c_out(c[1389]));
    fullAdder fa1296 (.a(s[1323]), .b(c[1322]), .c_in(c[1199]), .s(s[1390]), .c_out(c[1390]));
    fullAdder fa1297 (.a(s[1324]), .b(c[1323]), .c_in(c[1201]), .s(s[1391]), .c_out(c[1391]));
    fullAdder fa1298 (.a(s[1325]), .b(c[1324]), .c_in(c[1203]), .s(s[1392]), .c_out(c[1392]));
    fullAdder fa1299 (.a(s[1326]), .b(c[1325]), .c_in(c[1205]), .s(s[1393]), .c_out(c[1393]));
    fullAdder fa1300 (.a(s[1327]), .b(c[1326]), .c_in(c[1207]), .s(s[1394]), .c_out(c[1394]));
    fullAdder fa1301 (.a(s[1328]), .b(c[1327]), .c_in(c[1209]), .s(s[1395]), .c_out(c[1395]));
    fullAdder fa1302 (.a(s[1329]), .b(c[1328]), .c_in(c[1211]), .s(s[1396]), .c_out(c[1396]));
    fullAdder fa1303 (.a(s[1330]), .b(c[1329]), .c_in(s[1331]), .s(s[1397]), .c_out(c[1397]));
    fullAdder fa1304 (.a(s[1332]), .b(c[1330]), .c_in(c[445]), .s(s[1398]), .c_out(c[1398]));
    fullAdder fa1305 (.a(s[1333]), .b(c[1332]), .c_in(c[450]), .s(s[1399]), .c_out(c[1399]));
    fullAdder fa1306 (.a(s[1225]), .b(c[1341]), .c_in(c[1224]), .s(s[1400]), .c_out(c[1400]));
    fullAdder fa1307 (.a(s[1090]), .b(c[1342]), .c_in(c[1089]), .s(s[1401]), .c_out(c[1401]));
    // Stage 7 Reduction
    fullAdder fa1308 (.a(s[1242]), .b(c[1344]), .c_in(c[1241]), .s(s[1402]), .c_out(c[1402]));
    fullAdder fa1309 (.a(s[1246]), .b(c[1347]), .c_in(c[1245]), .s(s[1403]), .c_out(c[1403]));
    fullAdder fa1310 (.a(s[1356]), .b(c[1355]), .c_in(c[1256]), .s(s[1404]), .c_out(c[1404]));
    halfAdder ha96 (.a(s[1357]), .b(c[1356]), .s(s[1405]), .c_out(c[1405]));
    fullAdder fa1311 (.a(s[1358]), .b(c[1357]), .c_in(c[1259]), .s(s[1406]), .c_out(c[1406]));
    fullAdder fa1312 (.a(s[1359]), .b(c[1358]), .c_in(c[1261]), .s(s[1407]), .c_out(c[1407]));
    fullAdder fa1313 (.a(s[1360]), .b(c[1359]), .c_in(c[1263]), .s(s[1408]), .c_out(c[1408]));
    fullAdder fa1314 (.a(s[1361]), .b(c[1360]), .c_in(c[1265]), .s(s[1409]), .c_out(c[1409]));
    fullAdder fa1315 (.a(s[1362]), .b(c[1361]), .c_in(c[1267]), .s(s[1410]), .c_out(c[1410]));
    fullAdder fa1316 (.a(s[1363]), .b(c[1362]), .c_in(c[1269]), .s(s[1411]), .c_out(c[1411]));
    fullAdder fa1317 (.a(s[1364]), .b(c[1363]), .c_in(c[1271]), .s(s[1412]), .c_out(c[1412]));
    fullAdder fa1318 (.a(s[1365]), .b(c[1364]), .c_in(c[1273]), .s(s[1413]), .c_out(c[1413]));
    fullAdder fa1319 (.a(s[1366]), .b(c[1365]), .c_in(c[1275]), .s(s[1414]), .c_out(c[1414]));
    fullAdder fa1320 (.a(s[1367]), .b(c[1366]), .c_in(c[1277]), .s(s[1415]), .c_out(c[1415]));
    fullAdder fa1321 (.a(s[1368]), .b(c[1367]), .c_in(c[1279]), .s(s[1416]), .c_out(c[1416]));
    fullAdder fa1322 (.a(s[1369]), .b(c[1368]), .c_in(c[1281]), .s(s[1417]), .c_out(c[1417]));
    fullAdder fa1323 (.a(s[1370]), .b(c[1369]), .c_in(c[1283]), .s(s[1418]), .c_out(c[1418]));
    fullAdder fa1324 (.a(s[1371]), .b(c[1370]), .c_in(c[1285]), .s(s[1419]), .c_out(c[1419]));
    fullAdder fa1325 (.a(s[1372]), .b(c[1371]), .c_in(c[1287]), .s(s[1420]), .c_out(c[1420]));
    fullAdder fa1326 (.a(s[1373]), .b(c[1372]), .c_in(c[1289]), .s(s[1421]), .c_out(c[1421]));
    fullAdder fa1327 (.a(s[1374]), .b(c[1373]), .c_in(c[1291]), .s(s[1422]), .c_out(c[1422]));
    fullAdder fa1328 (.a(s[1375]), .b(c[1374]), .c_in(c[1293]), .s(s[1423]), .c_out(c[1423]));
    fullAdder fa1329 (.a(s[1376]), .b(c[1375]), .c_in(c[1295]), .s(s[1424]), .c_out(c[1424]));
    fullAdder fa1330 (.a(s[1377]), .b(c[1376]), .c_in(c[1297]), .s(s[1425]), .c_out(c[1425]));
    fullAdder fa1331 (.a(s[1378]), .b(c[1377]), .c_in(c[1299]), .s(s[1426]), .c_out(c[1426]));
    fullAdder fa1332 (.a(s[1379]), .b(c[1378]), .c_in(c[1301]), .s(s[1427]), .c_out(c[1427]));
    fullAdder fa1333 (.a(s[1380]), .b(c[1379]), .c_in(c[1303]), .s(s[1428]), .c_out(c[1428]));
    fullAdder fa1334 (.a(s[1381]), .b(c[1380]), .c_in(c[1305]), .s(s[1429]), .c_out(c[1429]));
    fullAdder fa1335 (.a(s[1382]), .b(c[1381]), .c_in(c[1307]), .s(s[1430]), .c_out(c[1430]));
    fullAdder fa1336 (.a(s[1383]), .b(c[1382]), .c_in(c[1309]), .s(s[1431]), .c_out(c[1431]));
    fullAdder fa1337 (.a(s[1384]), .b(c[1383]), .c_in(c[1311]), .s(s[1432]), .c_out(c[1432]));
    fullAdder fa1338 (.a(s[1385]), .b(c[1384]), .c_in(c[1313]), .s(s[1433]), .c_out(c[1433]));
    fullAdder fa1339 (.a(s[1386]), .b(c[1385]), .c_in(c[1315]), .s(s[1434]), .c_out(c[1434]));
    fullAdder fa1340 (.a(s[1387]), .b(c[1386]), .c_in(c[1317]), .s(s[1435]), .c_out(c[1435]));
    fullAdder fa1341 (.a(s[1388]), .b(c[1387]), .c_in(c[1319]), .s(s[1436]), .c_out(c[1436]));
    fullAdder fa1342 (.a(s[1389]), .b(c[1388]), .c_in(c[1321]), .s(s[1437]), .c_out(c[1437]));
    halfAdder ha97 (.a(s[1390]), .b(c[1389]), .s(s[1438]), .c_out(c[1438]));
    halfAdder ha98 (.a(s[1391]), .b(c[1390]), .s(s[1439]), .c_out(c[1439]));
    halfAdder ha99 (.a(s[1392]), .b(c[1391]), .s(s[1440]), .c_out(c[1440]));
    halfAdder ha100 (.a(s[1393]), .b(c[1392]), .s(s[1441]), .c_out(c[1441]));
    halfAdder ha101 (.a(s[1394]), .b(c[1393]), .s(s[1442]), .c_out(c[1442]));
    halfAdder ha102 (.a(s[1395]), .b(c[1394]), .s(s[1443]), .c_out(c[1443]));
    halfAdder ha103 (.a(s[1396]), .b(c[1395]), .s(s[1444]), .c_out(c[1444]));
    halfAdder ha104 (.a(s[1397]), .b(c[1396]), .s(s[1445]), .c_out(c[1445]));
    fullAdder fa1343 (.a(s[1398]), .b(c[1397]), .c_in(c[1331]), .s(s[1446]), .c_out(c[1446]));
    halfAdder ha105 (.a(s[1399]), .b(c[1398]), .s(s[1447]), .c_out(c[1447]));
    fullAdder fa1344 (.a(s[1334]), .b(c[1399]), .c_in(c[1333]), .s(s[1448]), .c_out(c[1448]));
    halfAdder ha106 (.a(s[1335]), .b(c[1334]), .s(s[1449]), .c_out(c[1449]));
    halfAdder ha107 (.a(s[1336]), .b(c[1335]), .s(s[1450]), .c_out(c[1450]));
    halfAdder ha108 (.a(s[1337]), .b(c[1336]), .s(s[1451]), .c_out(c[1451]));
    halfAdder ha109 (.a(s[1338]), .b(c[1337]), .s(s[1452]), .c_out(c[1452]));
    halfAdder ha110 (.a(s[1339]), .b(c[1338]), .s(s[1453]), .c_out(c[1453]));
    halfAdder ha111 (.a(s[1340]), .b(c[1339]), .s(s[1454]), .c_out(c[1454]));
    halfAdder ha112 (.a(s[1341]), .b(c[1340]), .s(s[1455]), .c_out(c[1455]));
    fullAdder fa1345 (.a(s[1226]), .b(c[1400]), .c_in(c[1225]), .s(s[1456]), .c_out(c[1456]));
    halfAdder ha113 (.a(s[1227]), .b(c[1226]), .s(s[1457]), .c_out(c[1457]));
    halfAdder ha114 (.a(s[1228]), .b(c[1227]), .s(s[1458]), .c_out(c[1458]));
    halfAdder ha115 (.a(s[1229]), .b(c[1228]), .s(s[1459]), .c_out(c[1459]));
    halfAdder ha116 (.a(s[1230]), .b(c[1229]), .s(s[1460]), .c_out(c[1460]));
    fullAdder fa1346 (.a(s[1091]), .b(c[1401]), .c_in(c[1090]), .s(s[1461]), .c_out(c[1461]));
    halfAdder ha117 (.a(s[1092]), .b(c[1091]), .s(s[1462]), .c_out(c[1462]));

endmodule